# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SRAM
#       Words            : 16384
#       Bits             : 32
#       Byte-Write       : 1
#       Aspect Ratio     : 4
#       Output Loading   : 1.3  (pf)
#       Data Slew        : 2.0  (ns)
#       CK Slew          : 2.0  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2018/01/11 13:38:03
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SRAM
CLASS BLOCK ;
FOREIGN SRAM 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 1920.140 BY 1391.600 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 1919.020 1380.180 1920.140 1383.420 ;
  LAYER metal3 ;
  RECT 1919.020 1380.180 1920.140 1383.420 ;
  LAYER metal2 ;
  RECT 1919.020 1380.180 1920.140 1383.420 ;
  LAYER metal1 ;
  RECT 1919.020 1380.180 1920.140 1383.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1372.340 1920.140 1375.580 ;
  LAYER metal3 ;
  RECT 1919.020 1372.340 1920.140 1375.580 ;
  LAYER metal2 ;
  RECT 1919.020 1372.340 1920.140 1375.580 ;
  LAYER metal1 ;
  RECT 1919.020 1372.340 1920.140 1375.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1364.500 1920.140 1367.740 ;
  LAYER metal3 ;
  RECT 1919.020 1364.500 1920.140 1367.740 ;
  LAYER metal2 ;
  RECT 1919.020 1364.500 1920.140 1367.740 ;
  LAYER metal1 ;
  RECT 1919.020 1364.500 1920.140 1367.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1356.660 1920.140 1359.900 ;
  LAYER metal3 ;
  RECT 1919.020 1356.660 1920.140 1359.900 ;
  LAYER metal2 ;
  RECT 1919.020 1356.660 1920.140 1359.900 ;
  LAYER metal1 ;
  RECT 1919.020 1356.660 1920.140 1359.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1348.820 1920.140 1352.060 ;
  LAYER metal3 ;
  RECT 1919.020 1348.820 1920.140 1352.060 ;
  LAYER metal2 ;
  RECT 1919.020 1348.820 1920.140 1352.060 ;
  LAYER metal1 ;
  RECT 1919.020 1348.820 1920.140 1352.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1340.980 1920.140 1344.220 ;
  LAYER metal3 ;
  RECT 1919.020 1340.980 1920.140 1344.220 ;
  LAYER metal2 ;
  RECT 1919.020 1340.980 1920.140 1344.220 ;
  LAYER metal1 ;
  RECT 1919.020 1340.980 1920.140 1344.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1301.780 1920.140 1305.020 ;
  LAYER metal3 ;
  RECT 1919.020 1301.780 1920.140 1305.020 ;
  LAYER metal2 ;
  RECT 1919.020 1301.780 1920.140 1305.020 ;
  LAYER metal1 ;
  RECT 1919.020 1301.780 1920.140 1305.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1293.940 1920.140 1297.180 ;
  LAYER metal3 ;
  RECT 1919.020 1293.940 1920.140 1297.180 ;
  LAYER metal2 ;
  RECT 1919.020 1293.940 1920.140 1297.180 ;
  LAYER metal1 ;
  RECT 1919.020 1293.940 1920.140 1297.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1286.100 1920.140 1289.340 ;
  LAYER metal3 ;
  RECT 1919.020 1286.100 1920.140 1289.340 ;
  LAYER metal2 ;
  RECT 1919.020 1286.100 1920.140 1289.340 ;
  LAYER metal1 ;
  RECT 1919.020 1286.100 1920.140 1289.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1278.260 1920.140 1281.500 ;
  LAYER metal3 ;
  RECT 1919.020 1278.260 1920.140 1281.500 ;
  LAYER metal2 ;
  RECT 1919.020 1278.260 1920.140 1281.500 ;
  LAYER metal1 ;
  RECT 1919.020 1278.260 1920.140 1281.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1270.420 1920.140 1273.660 ;
  LAYER metal3 ;
  RECT 1919.020 1270.420 1920.140 1273.660 ;
  LAYER metal2 ;
  RECT 1919.020 1270.420 1920.140 1273.660 ;
  LAYER metal1 ;
  RECT 1919.020 1270.420 1920.140 1273.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1262.580 1920.140 1265.820 ;
  LAYER metal3 ;
  RECT 1919.020 1262.580 1920.140 1265.820 ;
  LAYER metal2 ;
  RECT 1919.020 1262.580 1920.140 1265.820 ;
  LAYER metal1 ;
  RECT 1919.020 1262.580 1920.140 1265.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1223.380 1920.140 1226.620 ;
  LAYER metal3 ;
  RECT 1919.020 1223.380 1920.140 1226.620 ;
  LAYER metal2 ;
  RECT 1919.020 1223.380 1920.140 1226.620 ;
  LAYER metal1 ;
  RECT 1919.020 1223.380 1920.140 1226.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1215.540 1920.140 1218.780 ;
  LAYER metal3 ;
  RECT 1919.020 1215.540 1920.140 1218.780 ;
  LAYER metal2 ;
  RECT 1919.020 1215.540 1920.140 1218.780 ;
  LAYER metal1 ;
  RECT 1919.020 1215.540 1920.140 1218.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1207.700 1920.140 1210.940 ;
  LAYER metal3 ;
  RECT 1919.020 1207.700 1920.140 1210.940 ;
  LAYER metal2 ;
  RECT 1919.020 1207.700 1920.140 1210.940 ;
  LAYER metal1 ;
  RECT 1919.020 1207.700 1920.140 1210.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1199.860 1920.140 1203.100 ;
  LAYER metal3 ;
  RECT 1919.020 1199.860 1920.140 1203.100 ;
  LAYER metal2 ;
  RECT 1919.020 1199.860 1920.140 1203.100 ;
  LAYER metal1 ;
  RECT 1919.020 1199.860 1920.140 1203.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1192.020 1920.140 1195.260 ;
  LAYER metal3 ;
  RECT 1919.020 1192.020 1920.140 1195.260 ;
  LAYER metal2 ;
  RECT 1919.020 1192.020 1920.140 1195.260 ;
  LAYER metal1 ;
  RECT 1919.020 1192.020 1920.140 1195.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1184.180 1920.140 1187.420 ;
  LAYER metal3 ;
  RECT 1919.020 1184.180 1920.140 1187.420 ;
  LAYER metal2 ;
  RECT 1919.020 1184.180 1920.140 1187.420 ;
  LAYER metal1 ;
  RECT 1919.020 1184.180 1920.140 1187.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1144.980 1920.140 1148.220 ;
  LAYER metal3 ;
  RECT 1919.020 1144.980 1920.140 1148.220 ;
  LAYER metal2 ;
  RECT 1919.020 1144.980 1920.140 1148.220 ;
  LAYER metal1 ;
  RECT 1919.020 1144.980 1920.140 1148.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1137.140 1920.140 1140.380 ;
  LAYER metal3 ;
  RECT 1919.020 1137.140 1920.140 1140.380 ;
  LAYER metal2 ;
  RECT 1919.020 1137.140 1920.140 1140.380 ;
  LAYER metal1 ;
  RECT 1919.020 1137.140 1920.140 1140.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1129.300 1920.140 1132.540 ;
  LAYER metal3 ;
  RECT 1919.020 1129.300 1920.140 1132.540 ;
  LAYER metal2 ;
  RECT 1919.020 1129.300 1920.140 1132.540 ;
  LAYER metal1 ;
  RECT 1919.020 1129.300 1920.140 1132.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1121.460 1920.140 1124.700 ;
  LAYER metal3 ;
  RECT 1919.020 1121.460 1920.140 1124.700 ;
  LAYER metal2 ;
  RECT 1919.020 1121.460 1920.140 1124.700 ;
  LAYER metal1 ;
  RECT 1919.020 1121.460 1920.140 1124.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1113.620 1920.140 1116.860 ;
  LAYER metal3 ;
  RECT 1919.020 1113.620 1920.140 1116.860 ;
  LAYER metal2 ;
  RECT 1919.020 1113.620 1920.140 1116.860 ;
  LAYER metal1 ;
  RECT 1919.020 1113.620 1920.140 1116.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1105.780 1920.140 1109.020 ;
  LAYER metal3 ;
  RECT 1919.020 1105.780 1920.140 1109.020 ;
  LAYER metal2 ;
  RECT 1919.020 1105.780 1920.140 1109.020 ;
  LAYER metal1 ;
  RECT 1919.020 1105.780 1920.140 1109.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1066.580 1920.140 1069.820 ;
  LAYER metal3 ;
  RECT 1919.020 1066.580 1920.140 1069.820 ;
  LAYER metal2 ;
  RECT 1919.020 1066.580 1920.140 1069.820 ;
  LAYER metal1 ;
  RECT 1919.020 1066.580 1920.140 1069.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1058.740 1920.140 1061.980 ;
  LAYER metal3 ;
  RECT 1919.020 1058.740 1920.140 1061.980 ;
  LAYER metal2 ;
  RECT 1919.020 1058.740 1920.140 1061.980 ;
  LAYER metal1 ;
  RECT 1919.020 1058.740 1920.140 1061.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1050.900 1920.140 1054.140 ;
  LAYER metal3 ;
  RECT 1919.020 1050.900 1920.140 1054.140 ;
  LAYER metal2 ;
  RECT 1919.020 1050.900 1920.140 1054.140 ;
  LAYER metal1 ;
  RECT 1919.020 1050.900 1920.140 1054.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1043.060 1920.140 1046.300 ;
  LAYER metal3 ;
  RECT 1919.020 1043.060 1920.140 1046.300 ;
  LAYER metal2 ;
  RECT 1919.020 1043.060 1920.140 1046.300 ;
  LAYER metal1 ;
  RECT 1919.020 1043.060 1920.140 1046.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1035.220 1920.140 1038.460 ;
  LAYER metal3 ;
  RECT 1919.020 1035.220 1920.140 1038.460 ;
  LAYER metal2 ;
  RECT 1919.020 1035.220 1920.140 1038.460 ;
  LAYER metal1 ;
  RECT 1919.020 1035.220 1920.140 1038.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1027.380 1920.140 1030.620 ;
  LAYER metal3 ;
  RECT 1919.020 1027.380 1920.140 1030.620 ;
  LAYER metal2 ;
  RECT 1919.020 1027.380 1920.140 1030.620 ;
  LAYER metal1 ;
  RECT 1919.020 1027.380 1920.140 1030.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 988.180 1920.140 991.420 ;
  LAYER metal3 ;
  RECT 1919.020 988.180 1920.140 991.420 ;
  LAYER metal2 ;
  RECT 1919.020 988.180 1920.140 991.420 ;
  LAYER metal1 ;
  RECT 1919.020 988.180 1920.140 991.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 980.340 1920.140 983.580 ;
  LAYER metal3 ;
  RECT 1919.020 980.340 1920.140 983.580 ;
  LAYER metal2 ;
  RECT 1919.020 980.340 1920.140 983.580 ;
  LAYER metal1 ;
  RECT 1919.020 980.340 1920.140 983.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 972.500 1920.140 975.740 ;
  LAYER metal3 ;
  RECT 1919.020 972.500 1920.140 975.740 ;
  LAYER metal2 ;
  RECT 1919.020 972.500 1920.140 975.740 ;
  LAYER metal1 ;
  RECT 1919.020 972.500 1920.140 975.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 964.660 1920.140 967.900 ;
  LAYER metal3 ;
  RECT 1919.020 964.660 1920.140 967.900 ;
  LAYER metal2 ;
  RECT 1919.020 964.660 1920.140 967.900 ;
  LAYER metal1 ;
  RECT 1919.020 964.660 1920.140 967.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 956.820 1920.140 960.060 ;
  LAYER metal3 ;
  RECT 1919.020 956.820 1920.140 960.060 ;
  LAYER metal2 ;
  RECT 1919.020 956.820 1920.140 960.060 ;
  LAYER metal1 ;
  RECT 1919.020 956.820 1920.140 960.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 948.980 1920.140 952.220 ;
  LAYER metal3 ;
  RECT 1919.020 948.980 1920.140 952.220 ;
  LAYER metal2 ;
  RECT 1919.020 948.980 1920.140 952.220 ;
  LAYER metal1 ;
  RECT 1919.020 948.980 1920.140 952.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 909.780 1920.140 913.020 ;
  LAYER metal3 ;
  RECT 1919.020 909.780 1920.140 913.020 ;
  LAYER metal2 ;
  RECT 1919.020 909.780 1920.140 913.020 ;
  LAYER metal1 ;
  RECT 1919.020 909.780 1920.140 913.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 901.940 1920.140 905.180 ;
  LAYER metal3 ;
  RECT 1919.020 901.940 1920.140 905.180 ;
  LAYER metal2 ;
  RECT 1919.020 901.940 1920.140 905.180 ;
  LAYER metal1 ;
  RECT 1919.020 901.940 1920.140 905.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 894.100 1920.140 897.340 ;
  LAYER metal3 ;
  RECT 1919.020 894.100 1920.140 897.340 ;
  LAYER metal2 ;
  RECT 1919.020 894.100 1920.140 897.340 ;
  LAYER metal1 ;
  RECT 1919.020 894.100 1920.140 897.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 886.260 1920.140 889.500 ;
  LAYER metal3 ;
  RECT 1919.020 886.260 1920.140 889.500 ;
  LAYER metal2 ;
  RECT 1919.020 886.260 1920.140 889.500 ;
  LAYER metal1 ;
  RECT 1919.020 886.260 1920.140 889.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 878.420 1920.140 881.660 ;
  LAYER metal3 ;
  RECT 1919.020 878.420 1920.140 881.660 ;
  LAYER metal2 ;
  RECT 1919.020 878.420 1920.140 881.660 ;
  LAYER metal1 ;
  RECT 1919.020 878.420 1920.140 881.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 870.580 1920.140 873.820 ;
  LAYER metal3 ;
  RECT 1919.020 870.580 1920.140 873.820 ;
  LAYER metal2 ;
  RECT 1919.020 870.580 1920.140 873.820 ;
  LAYER metal1 ;
  RECT 1919.020 870.580 1920.140 873.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 831.380 1920.140 834.620 ;
  LAYER metal3 ;
  RECT 1919.020 831.380 1920.140 834.620 ;
  LAYER metal2 ;
  RECT 1919.020 831.380 1920.140 834.620 ;
  LAYER metal1 ;
  RECT 1919.020 831.380 1920.140 834.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 823.540 1920.140 826.780 ;
  LAYER metal3 ;
  RECT 1919.020 823.540 1920.140 826.780 ;
  LAYER metal2 ;
  RECT 1919.020 823.540 1920.140 826.780 ;
  LAYER metal1 ;
  RECT 1919.020 823.540 1920.140 826.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 815.700 1920.140 818.940 ;
  LAYER metal3 ;
  RECT 1919.020 815.700 1920.140 818.940 ;
  LAYER metal2 ;
  RECT 1919.020 815.700 1920.140 818.940 ;
  LAYER metal1 ;
  RECT 1919.020 815.700 1920.140 818.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 807.860 1920.140 811.100 ;
  LAYER metal3 ;
  RECT 1919.020 807.860 1920.140 811.100 ;
  LAYER metal2 ;
  RECT 1919.020 807.860 1920.140 811.100 ;
  LAYER metal1 ;
  RECT 1919.020 807.860 1920.140 811.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 800.020 1920.140 803.260 ;
  LAYER metal3 ;
  RECT 1919.020 800.020 1920.140 803.260 ;
  LAYER metal2 ;
  RECT 1919.020 800.020 1920.140 803.260 ;
  LAYER metal1 ;
  RECT 1919.020 800.020 1920.140 803.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 792.180 1920.140 795.420 ;
  LAYER metal3 ;
  RECT 1919.020 792.180 1920.140 795.420 ;
  LAYER metal2 ;
  RECT 1919.020 792.180 1920.140 795.420 ;
  LAYER metal1 ;
  RECT 1919.020 792.180 1920.140 795.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 752.980 1920.140 756.220 ;
  LAYER metal3 ;
  RECT 1919.020 752.980 1920.140 756.220 ;
  LAYER metal2 ;
  RECT 1919.020 752.980 1920.140 756.220 ;
  LAYER metal1 ;
  RECT 1919.020 752.980 1920.140 756.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 745.140 1920.140 748.380 ;
  LAYER metal3 ;
  RECT 1919.020 745.140 1920.140 748.380 ;
  LAYER metal2 ;
  RECT 1919.020 745.140 1920.140 748.380 ;
  LAYER metal1 ;
  RECT 1919.020 745.140 1920.140 748.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 737.300 1920.140 740.540 ;
  LAYER metal3 ;
  RECT 1919.020 737.300 1920.140 740.540 ;
  LAYER metal2 ;
  RECT 1919.020 737.300 1920.140 740.540 ;
  LAYER metal1 ;
  RECT 1919.020 737.300 1920.140 740.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 729.460 1920.140 732.700 ;
  LAYER metal3 ;
  RECT 1919.020 729.460 1920.140 732.700 ;
  LAYER metal2 ;
  RECT 1919.020 729.460 1920.140 732.700 ;
  LAYER metal1 ;
  RECT 1919.020 729.460 1920.140 732.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 721.620 1920.140 724.860 ;
  LAYER metal3 ;
  RECT 1919.020 721.620 1920.140 724.860 ;
  LAYER metal2 ;
  RECT 1919.020 721.620 1920.140 724.860 ;
  LAYER metal1 ;
  RECT 1919.020 721.620 1920.140 724.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 713.780 1920.140 717.020 ;
  LAYER metal3 ;
  RECT 1919.020 713.780 1920.140 717.020 ;
  LAYER metal2 ;
  RECT 1919.020 713.780 1920.140 717.020 ;
  LAYER metal1 ;
  RECT 1919.020 713.780 1920.140 717.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 674.580 1920.140 677.820 ;
  LAYER metal3 ;
  RECT 1919.020 674.580 1920.140 677.820 ;
  LAYER metal2 ;
  RECT 1919.020 674.580 1920.140 677.820 ;
  LAYER metal1 ;
  RECT 1919.020 674.580 1920.140 677.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 666.740 1920.140 669.980 ;
  LAYER metal3 ;
  RECT 1919.020 666.740 1920.140 669.980 ;
  LAYER metal2 ;
  RECT 1919.020 666.740 1920.140 669.980 ;
  LAYER metal1 ;
  RECT 1919.020 666.740 1920.140 669.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 658.900 1920.140 662.140 ;
  LAYER metal3 ;
  RECT 1919.020 658.900 1920.140 662.140 ;
  LAYER metal2 ;
  RECT 1919.020 658.900 1920.140 662.140 ;
  LAYER metal1 ;
  RECT 1919.020 658.900 1920.140 662.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 651.060 1920.140 654.300 ;
  LAYER metal3 ;
  RECT 1919.020 651.060 1920.140 654.300 ;
  LAYER metal2 ;
  RECT 1919.020 651.060 1920.140 654.300 ;
  LAYER metal1 ;
  RECT 1919.020 651.060 1920.140 654.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 643.220 1920.140 646.460 ;
  LAYER metal3 ;
  RECT 1919.020 643.220 1920.140 646.460 ;
  LAYER metal2 ;
  RECT 1919.020 643.220 1920.140 646.460 ;
  LAYER metal1 ;
  RECT 1919.020 643.220 1920.140 646.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 635.380 1920.140 638.620 ;
  LAYER metal3 ;
  RECT 1919.020 635.380 1920.140 638.620 ;
  LAYER metal2 ;
  RECT 1919.020 635.380 1920.140 638.620 ;
  LAYER metal1 ;
  RECT 1919.020 635.380 1920.140 638.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 596.180 1920.140 599.420 ;
  LAYER metal3 ;
  RECT 1919.020 596.180 1920.140 599.420 ;
  LAYER metal2 ;
  RECT 1919.020 596.180 1920.140 599.420 ;
  LAYER metal1 ;
  RECT 1919.020 596.180 1920.140 599.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 588.340 1920.140 591.580 ;
  LAYER metal3 ;
  RECT 1919.020 588.340 1920.140 591.580 ;
  LAYER metal2 ;
  RECT 1919.020 588.340 1920.140 591.580 ;
  LAYER metal1 ;
  RECT 1919.020 588.340 1920.140 591.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 580.500 1920.140 583.740 ;
  LAYER metal3 ;
  RECT 1919.020 580.500 1920.140 583.740 ;
  LAYER metal2 ;
  RECT 1919.020 580.500 1920.140 583.740 ;
  LAYER metal1 ;
  RECT 1919.020 580.500 1920.140 583.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 572.660 1920.140 575.900 ;
  LAYER metal3 ;
  RECT 1919.020 572.660 1920.140 575.900 ;
  LAYER metal2 ;
  RECT 1919.020 572.660 1920.140 575.900 ;
  LAYER metal1 ;
  RECT 1919.020 572.660 1920.140 575.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 564.820 1920.140 568.060 ;
  LAYER metal3 ;
  RECT 1919.020 564.820 1920.140 568.060 ;
  LAYER metal2 ;
  RECT 1919.020 564.820 1920.140 568.060 ;
  LAYER metal1 ;
  RECT 1919.020 564.820 1920.140 568.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 556.980 1920.140 560.220 ;
  LAYER metal3 ;
  RECT 1919.020 556.980 1920.140 560.220 ;
  LAYER metal2 ;
  RECT 1919.020 556.980 1920.140 560.220 ;
  LAYER metal1 ;
  RECT 1919.020 556.980 1920.140 560.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 517.780 1920.140 521.020 ;
  LAYER metal3 ;
  RECT 1919.020 517.780 1920.140 521.020 ;
  LAYER metal2 ;
  RECT 1919.020 517.780 1920.140 521.020 ;
  LAYER metal1 ;
  RECT 1919.020 517.780 1920.140 521.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 509.940 1920.140 513.180 ;
  LAYER metal3 ;
  RECT 1919.020 509.940 1920.140 513.180 ;
  LAYER metal2 ;
  RECT 1919.020 509.940 1920.140 513.180 ;
  LAYER metal1 ;
  RECT 1919.020 509.940 1920.140 513.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 502.100 1920.140 505.340 ;
  LAYER metal3 ;
  RECT 1919.020 502.100 1920.140 505.340 ;
  LAYER metal2 ;
  RECT 1919.020 502.100 1920.140 505.340 ;
  LAYER metal1 ;
  RECT 1919.020 502.100 1920.140 505.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 494.260 1920.140 497.500 ;
  LAYER metal3 ;
  RECT 1919.020 494.260 1920.140 497.500 ;
  LAYER metal2 ;
  RECT 1919.020 494.260 1920.140 497.500 ;
  LAYER metal1 ;
  RECT 1919.020 494.260 1920.140 497.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 486.420 1920.140 489.660 ;
  LAYER metal3 ;
  RECT 1919.020 486.420 1920.140 489.660 ;
  LAYER metal2 ;
  RECT 1919.020 486.420 1920.140 489.660 ;
  LAYER metal1 ;
  RECT 1919.020 486.420 1920.140 489.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 478.580 1920.140 481.820 ;
  LAYER metal3 ;
  RECT 1919.020 478.580 1920.140 481.820 ;
  LAYER metal2 ;
  RECT 1919.020 478.580 1920.140 481.820 ;
  LAYER metal1 ;
  RECT 1919.020 478.580 1920.140 481.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 439.380 1920.140 442.620 ;
  LAYER metal3 ;
  RECT 1919.020 439.380 1920.140 442.620 ;
  LAYER metal2 ;
  RECT 1919.020 439.380 1920.140 442.620 ;
  LAYER metal1 ;
  RECT 1919.020 439.380 1920.140 442.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 431.540 1920.140 434.780 ;
  LAYER metal3 ;
  RECT 1919.020 431.540 1920.140 434.780 ;
  LAYER metal2 ;
  RECT 1919.020 431.540 1920.140 434.780 ;
  LAYER metal1 ;
  RECT 1919.020 431.540 1920.140 434.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 423.700 1920.140 426.940 ;
  LAYER metal3 ;
  RECT 1919.020 423.700 1920.140 426.940 ;
  LAYER metal2 ;
  RECT 1919.020 423.700 1920.140 426.940 ;
  LAYER metal1 ;
  RECT 1919.020 423.700 1920.140 426.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 415.860 1920.140 419.100 ;
  LAYER metal3 ;
  RECT 1919.020 415.860 1920.140 419.100 ;
  LAYER metal2 ;
  RECT 1919.020 415.860 1920.140 419.100 ;
  LAYER metal1 ;
  RECT 1919.020 415.860 1920.140 419.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 408.020 1920.140 411.260 ;
  LAYER metal3 ;
  RECT 1919.020 408.020 1920.140 411.260 ;
  LAYER metal2 ;
  RECT 1919.020 408.020 1920.140 411.260 ;
  LAYER metal1 ;
  RECT 1919.020 408.020 1920.140 411.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 400.180 1920.140 403.420 ;
  LAYER metal3 ;
  RECT 1919.020 400.180 1920.140 403.420 ;
  LAYER metal2 ;
  RECT 1919.020 400.180 1920.140 403.420 ;
  LAYER metal1 ;
  RECT 1919.020 400.180 1920.140 403.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 360.980 1920.140 364.220 ;
  LAYER metal3 ;
  RECT 1919.020 360.980 1920.140 364.220 ;
  LAYER metal2 ;
  RECT 1919.020 360.980 1920.140 364.220 ;
  LAYER metal1 ;
  RECT 1919.020 360.980 1920.140 364.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 353.140 1920.140 356.380 ;
  LAYER metal3 ;
  RECT 1919.020 353.140 1920.140 356.380 ;
  LAYER metal2 ;
  RECT 1919.020 353.140 1920.140 356.380 ;
  LAYER metal1 ;
  RECT 1919.020 353.140 1920.140 356.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 345.300 1920.140 348.540 ;
  LAYER metal3 ;
  RECT 1919.020 345.300 1920.140 348.540 ;
  LAYER metal2 ;
  RECT 1919.020 345.300 1920.140 348.540 ;
  LAYER metal1 ;
  RECT 1919.020 345.300 1920.140 348.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 337.460 1920.140 340.700 ;
  LAYER metal3 ;
  RECT 1919.020 337.460 1920.140 340.700 ;
  LAYER metal2 ;
  RECT 1919.020 337.460 1920.140 340.700 ;
  LAYER metal1 ;
  RECT 1919.020 337.460 1920.140 340.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 329.620 1920.140 332.860 ;
  LAYER metal3 ;
  RECT 1919.020 329.620 1920.140 332.860 ;
  LAYER metal2 ;
  RECT 1919.020 329.620 1920.140 332.860 ;
  LAYER metal1 ;
  RECT 1919.020 329.620 1920.140 332.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 321.780 1920.140 325.020 ;
  LAYER metal3 ;
  RECT 1919.020 321.780 1920.140 325.020 ;
  LAYER metal2 ;
  RECT 1919.020 321.780 1920.140 325.020 ;
  LAYER metal1 ;
  RECT 1919.020 321.780 1920.140 325.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 282.580 1920.140 285.820 ;
  LAYER metal3 ;
  RECT 1919.020 282.580 1920.140 285.820 ;
  LAYER metal2 ;
  RECT 1919.020 282.580 1920.140 285.820 ;
  LAYER metal1 ;
  RECT 1919.020 282.580 1920.140 285.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 274.740 1920.140 277.980 ;
  LAYER metal3 ;
  RECT 1919.020 274.740 1920.140 277.980 ;
  LAYER metal2 ;
  RECT 1919.020 274.740 1920.140 277.980 ;
  LAYER metal1 ;
  RECT 1919.020 274.740 1920.140 277.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 266.900 1920.140 270.140 ;
  LAYER metal3 ;
  RECT 1919.020 266.900 1920.140 270.140 ;
  LAYER metal2 ;
  RECT 1919.020 266.900 1920.140 270.140 ;
  LAYER metal1 ;
  RECT 1919.020 266.900 1920.140 270.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 259.060 1920.140 262.300 ;
  LAYER metal3 ;
  RECT 1919.020 259.060 1920.140 262.300 ;
  LAYER metal2 ;
  RECT 1919.020 259.060 1920.140 262.300 ;
  LAYER metal1 ;
  RECT 1919.020 259.060 1920.140 262.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 251.220 1920.140 254.460 ;
  LAYER metal3 ;
  RECT 1919.020 251.220 1920.140 254.460 ;
  LAYER metal2 ;
  RECT 1919.020 251.220 1920.140 254.460 ;
  LAYER metal1 ;
  RECT 1919.020 251.220 1920.140 254.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 243.380 1920.140 246.620 ;
  LAYER metal3 ;
  RECT 1919.020 243.380 1920.140 246.620 ;
  LAYER metal2 ;
  RECT 1919.020 243.380 1920.140 246.620 ;
  LAYER metal1 ;
  RECT 1919.020 243.380 1920.140 246.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 204.180 1920.140 207.420 ;
  LAYER metal3 ;
  RECT 1919.020 204.180 1920.140 207.420 ;
  LAYER metal2 ;
  RECT 1919.020 204.180 1920.140 207.420 ;
  LAYER metal1 ;
  RECT 1919.020 204.180 1920.140 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 196.340 1920.140 199.580 ;
  LAYER metal3 ;
  RECT 1919.020 196.340 1920.140 199.580 ;
  LAYER metal2 ;
  RECT 1919.020 196.340 1920.140 199.580 ;
  LAYER metal1 ;
  RECT 1919.020 196.340 1920.140 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 188.500 1920.140 191.740 ;
  LAYER metal3 ;
  RECT 1919.020 188.500 1920.140 191.740 ;
  LAYER metal2 ;
  RECT 1919.020 188.500 1920.140 191.740 ;
  LAYER metal1 ;
  RECT 1919.020 188.500 1920.140 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 180.660 1920.140 183.900 ;
  LAYER metal3 ;
  RECT 1919.020 180.660 1920.140 183.900 ;
  LAYER metal2 ;
  RECT 1919.020 180.660 1920.140 183.900 ;
  LAYER metal1 ;
  RECT 1919.020 180.660 1920.140 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 172.820 1920.140 176.060 ;
  LAYER metal3 ;
  RECT 1919.020 172.820 1920.140 176.060 ;
  LAYER metal2 ;
  RECT 1919.020 172.820 1920.140 176.060 ;
  LAYER metal1 ;
  RECT 1919.020 172.820 1920.140 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 164.980 1920.140 168.220 ;
  LAYER metal3 ;
  RECT 1919.020 164.980 1920.140 168.220 ;
  LAYER metal2 ;
  RECT 1919.020 164.980 1920.140 168.220 ;
  LAYER metal1 ;
  RECT 1919.020 164.980 1920.140 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 125.780 1920.140 129.020 ;
  LAYER metal3 ;
  RECT 1919.020 125.780 1920.140 129.020 ;
  LAYER metal2 ;
  RECT 1919.020 125.780 1920.140 129.020 ;
  LAYER metal1 ;
  RECT 1919.020 125.780 1920.140 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 117.940 1920.140 121.180 ;
  LAYER metal3 ;
  RECT 1919.020 117.940 1920.140 121.180 ;
  LAYER metal2 ;
  RECT 1919.020 117.940 1920.140 121.180 ;
  LAYER metal1 ;
  RECT 1919.020 117.940 1920.140 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 110.100 1920.140 113.340 ;
  LAYER metal3 ;
  RECT 1919.020 110.100 1920.140 113.340 ;
  LAYER metal2 ;
  RECT 1919.020 110.100 1920.140 113.340 ;
  LAYER metal1 ;
  RECT 1919.020 110.100 1920.140 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 102.260 1920.140 105.500 ;
  LAYER metal3 ;
  RECT 1919.020 102.260 1920.140 105.500 ;
  LAYER metal2 ;
  RECT 1919.020 102.260 1920.140 105.500 ;
  LAYER metal1 ;
  RECT 1919.020 102.260 1920.140 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 94.420 1920.140 97.660 ;
  LAYER metal3 ;
  RECT 1919.020 94.420 1920.140 97.660 ;
  LAYER metal2 ;
  RECT 1919.020 94.420 1920.140 97.660 ;
  LAYER metal1 ;
  RECT 1919.020 94.420 1920.140 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 86.580 1920.140 89.820 ;
  LAYER metal3 ;
  RECT 1919.020 86.580 1920.140 89.820 ;
  LAYER metal2 ;
  RECT 1919.020 86.580 1920.140 89.820 ;
  LAYER metal1 ;
  RECT 1919.020 86.580 1920.140 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 47.380 1920.140 50.620 ;
  LAYER metal3 ;
  RECT 1919.020 47.380 1920.140 50.620 ;
  LAYER metal2 ;
  RECT 1919.020 47.380 1920.140 50.620 ;
  LAYER metal1 ;
  RECT 1919.020 47.380 1920.140 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 39.540 1920.140 42.780 ;
  LAYER metal3 ;
  RECT 1919.020 39.540 1920.140 42.780 ;
  LAYER metal2 ;
  RECT 1919.020 39.540 1920.140 42.780 ;
  LAYER metal1 ;
  RECT 1919.020 39.540 1920.140 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 31.700 1920.140 34.940 ;
  LAYER metal3 ;
  RECT 1919.020 31.700 1920.140 34.940 ;
  LAYER metal2 ;
  RECT 1919.020 31.700 1920.140 34.940 ;
  LAYER metal1 ;
  RECT 1919.020 31.700 1920.140 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 23.860 1920.140 27.100 ;
  LAYER metal3 ;
  RECT 1919.020 23.860 1920.140 27.100 ;
  LAYER metal2 ;
  RECT 1919.020 23.860 1920.140 27.100 ;
  LAYER metal1 ;
  RECT 1919.020 23.860 1920.140 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 16.020 1920.140 19.260 ;
  LAYER metal3 ;
  RECT 1919.020 16.020 1920.140 19.260 ;
  LAYER metal2 ;
  RECT 1919.020 16.020 1920.140 19.260 ;
  LAYER metal1 ;
  RECT 1919.020 16.020 1920.140 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 8.180 1920.140 11.420 ;
  LAYER metal3 ;
  RECT 1919.020 8.180 1920.140 11.420 ;
  LAYER metal2 ;
  RECT 1919.020 8.180 1920.140 11.420 ;
  LAYER metal1 ;
  RECT 1919.020 8.180 1920.140 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1380.180 1.120 1383.420 ;
  LAYER metal3 ;
  RECT 0.000 1380.180 1.120 1383.420 ;
  LAYER metal2 ;
  RECT 0.000 1380.180 1.120 1383.420 ;
  LAYER metal1 ;
  RECT 0.000 1380.180 1.120 1383.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1372.340 1.120 1375.580 ;
  LAYER metal3 ;
  RECT 0.000 1372.340 1.120 1375.580 ;
  LAYER metal2 ;
  RECT 0.000 1372.340 1.120 1375.580 ;
  LAYER metal1 ;
  RECT 0.000 1372.340 1.120 1375.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1364.500 1.120 1367.740 ;
  LAYER metal3 ;
  RECT 0.000 1364.500 1.120 1367.740 ;
  LAYER metal2 ;
  RECT 0.000 1364.500 1.120 1367.740 ;
  LAYER metal1 ;
  RECT 0.000 1364.500 1.120 1367.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1356.660 1.120 1359.900 ;
  LAYER metal3 ;
  RECT 0.000 1356.660 1.120 1359.900 ;
  LAYER metal2 ;
  RECT 0.000 1356.660 1.120 1359.900 ;
  LAYER metal1 ;
  RECT 0.000 1356.660 1.120 1359.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1348.820 1.120 1352.060 ;
  LAYER metal3 ;
  RECT 0.000 1348.820 1.120 1352.060 ;
  LAYER metal2 ;
  RECT 0.000 1348.820 1.120 1352.060 ;
  LAYER metal1 ;
  RECT 0.000 1348.820 1.120 1352.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1340.980 1.120 1344.220 ;
  LAYER metal3 ;
  RECT 0.000 1340.980 1.120 1344.220 ;
  LAYER metal2 ;
  RECT 0.000 1340.980 1.120 1344.220 ;
  LAYER metal1 ;
  RECT 0.000 1340.980 1.120 1344.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1301.780 1.120 1305.020 ;
  LAYER metal3 ;
  RECT 0.000 1301.780 1.120 1305.020 ;
  LAYER metal2 ;
  RECT 0.000 1301.780 1.120 1305.020 ;
  LAYER metal1 ;
  RECT 0.000 1301.780 1.120 1305.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1293.940 1.120 1297.180 ;
  LAYER metal3 ;
  RECT 0.000 1293.940 1.120 1297.180 ;
  LAYER metal2 ;
  RECT 0.000 1293.940 1.120 1297.180 ;
  LAYER metal1 ;
  RECT 0.000 1293.940 1.120 1297.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1286.100 1.120 1289.340 ;
  LAYER metal3 ;
  RECT 0.000 1286.100 1.120 1289.340 ;
  LAYER metal2 ;
  RECT 0.000 1286.100 1.120 1289.340 ;
  LAYER metal1 ;
  RECT 0.000 1286.100 1.120 1289.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1278.260 1.120 1281.500 ;
  LAYER metal3 ;
  RECT 0.000 1278.260 1.120 1281.500 ;
  LAYER metal2 ;
  RECT 0.000 1278.260 1.120 1281.500 ;
  LAYER metal1 ;
  RECT 0.000 1278.260 1.120 1281.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1270.420 1.120 1273.660 ;
  LAYER metal3 ;
  RECT 0.000 1270.420 1.120 1273.660 ;
  LAYER metal2 ;
  RECT 0.000 1270.420 1.120 1273.660 ;
  LAYER metal1 ;
  RECT 0.000 1270.420 1.120 1273.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1262.580 1.120 1265.820 ;
  LAYER metal3 ;
  RECT 0.000 1262.580 1.120 1265.820 ;
  LAYER metal2 ;
  RECT 0.000 1262.580 1.120 1265.820 ;
  LAYER metal1 ;
  RECT 0.000 1262.580 1.120 1265.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1223.380 1.120 1226.620 ;
  LAYER metal3 ;
  RECT 0.000 1223.380 1.120 1226.620 ;
  LAYER metal2 ;
  RECT 0.000 1223.380 1.120 1226.620 ;
  LAYER metal1 ;
  RECT 0.000 1223.380 1.120 1226.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1215.540 1.120 1218.780 ;
  LAYER metal3 ;
  RECT 0.000 1215.540 1.120 1218.780 ;
  LAYER metal2 ;
  RECT 0.000 1215.540 1.120 1218.780 ;
  LAYER metal1 ;
  RECT 0.000 1215.540 1.120 1218.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1207.700 1.120 1210.940 ;
  LAYER metal3 ;
  RECT 0.000 1207.700 1.120 1210.940 ;
  LAYER metal2 ;
  RECT 0.000 1207.700 1.120 1210.940 ;
  LAYER metal1 ;
  RECT 0.000 1207.700 1.120 1210.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1199.860 1.120 1203.100 ;
  LAYER metal3 ;
  RECT 0.000 1199.860 1.120 1203.100 ;
  LAYER metal2 ;
  RECT 0.000 1199.860 1.120 1203.100 ;
  LAYER metal1 ;
  RECT 0.000 1199.860 1.120 1203.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1192.020 1.120 1195.260 ;
  LAYER metal3 ;
  RECT 0.000 1192.020 1.120 1195.260 ;
  LAYER metal2 ;
  RECT 0.000 1192.020 1.120 1195.260 ;
  LAYER metal1 ;
  RECT 0.000 1192.020 1.120 1195.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1184.180 1.120 1187.420 ;
  LAYER metal3 ;
  RECT 0.000 1184.180 1.120 1187.420 ;
  LAYER metal2 ;
  RECT 0.000 1184.180 1.120 1187.420 ;
  LAYER metal1 ;
  RECT 0.000 1184.180 1.120 1187.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1144.980 1.120 1148.220 ;
  LAYER metal3 ;
  RECT 0.000 1144.980 1.120 1148.220 ;
  LAYER metal2 ;
  RECT 0.000 1144.980 1.120 1148.220 ;
  LAYER metal1 ;
  RECT 0.000 1144.980 1.120 1148.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1137.140 1.120 1140.380 ;
  LAYER metal3 ;
  RECT 0.000 1137.140 1.120 1140.380 ;
  LAYER metal2 ;
  RECT 0.000 1137.140 1.120 1140.380 ;
  LAYER metal1 ;
  RECT 0.000 1137.140 1.120 1140.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1129.300 1.120 1132.540 ;
  LAYER metal3 ;
  RECT 0.000 1129.300 1.120 1132.540 ;
  LAYER metal2 ;
  RECT 0.000 1129.300 1.120 1132.540 ;
  LAYER metal1 ;
  RECT 0.000 1129.300 1.120 1132.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1121.460 1.120 1124.700 ;
  LAYER metal3 ;
  RECT 0.000 1121.460 1.120 1124.700 ;
  LAYER metal2 ;
  RECT 0.000 1121.460 1.120 1124.700 ;
  LAYER metal1 ;
  RECT 0.000 1121.460 1.120 1124.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1113.620 1.120 1116.860 ;
  LAYER metal3 ;
  RECT 0.000 1113.620 1.120 1116.860 ;
  LAYER metal2 ;
  RECT 0.000 1113.620 1.120 1116.860 ;
  LAYER metal1 ;
  RECT 0.000 1113.620 1.120 1116.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1105.780 1.120 1109.020 ;
  LAYER metal3 ;
  RECT 0.000 1105.780 1.120 1109.020 ;
  LAYER metal2 ;
  RECT 0.000 1105.780 1.120 1109.020 ;
  LAYER metal1 ;
  RECT 0.000 1105.780 1.120 1109.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1066.580 1.120 1069.820 ;
  LAYER metal3 ;
  RECT 0.000 1066.580 1.120 1069.820 ;
  LAYER metal2 ;
  RECT 0.000 1066.580 1.120 1069.820 ;
  LAYER metal1 ;
  RECT 0.000 1066.580 1.120 1069.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1058.740 1.120 1061.980 ;
  LAYER metal3 ;
  RECT 0.000 1058.740 1.120 1061.980 ;
  LAYER metal2 ;
  RECT 0.000 1058.740 1.120 1061.980 ;
  LAYER metal1 ;
  RECT 0.000 1058.740 1.120 1061.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1050.900 1.120 1054.140 ;
  LAYER metal3 ;
  RECT 0.000 1050.900 1.120 1054.140 ;
  LAYER metal2 ;
  RECT 0.000 1050.900 1.120 1054.140 ;
  LAYER metal1 ;
  RECT 0.000 1050.900 1.120 1054.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1043.060 1.120 1046.300 ;
  LAYER metal3 ;
  RECT 0.000 1043.060 1.120 1046.300 ;
  LAYER metal2 ;
  RECT 0.000 1043.060 1.120 1046.300 ;
  LAYER metal1 ;
  RECT 0.000 1043.060 1.120 1046.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1035.220 1.120 1038.460 ;
  LAYER metal3 ;
  RECT 0.000 1035.220 1.120 1038.460 ;
  LAYER metal2 ;
  RECT 0.000 1035.220 1.120 1038.460 ;
  LAYER metal1 ;
  RECT 0.000 1035.220 1.120 1038.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1027.380 1.120 1030.620 ;
  LAYER metal3 ;
  RECT 0.000 1027.380 1.120 1030.620 ;
  LAYER metal2 ;
  RECT 0.000 1027.380 1.120 1030.620 ;
  LAYER metal1 ;
  RECT 0.000 1027.380 1.120 1030.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 988.180 1.120 991.420 ;
  LAYER metal3 ;
  RECT 0.000 988.180 1.120 991.420 ;
  LAYER metal2 ;
  RECT 0.000 988.180 1.120 991.420 ;
  LAYER metal1 ;
  RECT 0.000 988.180 1.120 991.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 980.340 1.120 983.580 ;
  LAYER metal3 ;
  RECT 0.000 980.340 1.120 983.580 ;
  LAYER metal2 ;
  RECT 0.000 980.340 1.120 983.580 ;
  LAYER metal1 ;
  RECT 0.000 980.340 1.120 983.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 972.500 1.120 975.740 ;
  LAYER metal3 ;
  RECT 0.000 972.500 1.120 975.740 ;
  LAYER metal2 ;
  RECT 0.000 972.500 1.120 975.740 ;
  LAYER metal1 ;
  RECT 0.000 972.500 1.120 975.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 964.660 1.120 967.900 ;
  LAYER metal3 ;
  RECT 0.000 964.660 1.120 967.900 ;
  LAYER metal2 ;
  RECT 0.000 964.660 1.120 967.900 ;
  LAYER metal1 ;
  RECT 0.000 964.660 1.120 967.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 956.820 1.120 960.060 ;
  LAYER metal3 ;
  RECT 0.000 956.820 1.120 960.060 ;
  LAYER metal2 ;
  RECT 0.000 956.820 1.120 960.060 ;
  LAYER metal1 ;
  RECT 0.000 956.820 1.120 960.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 948.980 1.120 952.220 ;
  LAYER metal3 ;
  RECT 0.000 948.980 1.120 952.220 ;
  LAYER metal2 ;
  RECT 0.000 948.980 1.120 952.220 ;
  LAYER metal1 ;
  RECT 0.000 948.980 1.120 952.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 909.780 1.120 913.020 ;
  LAYER metal3 ;
  RECT 0.000 909.780 1.120 913.020 ;
  LAYER metal2 ;
  RECT 0.000 909.780 1.120 913.020 ;
  LAYER metal1 ;
  RECT 0.000 909.780 1.120 913.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 901.940 1.120 905.180 ;
  LAYER metal3 ;
  RECT 0.000 901.940 1.120 905.180 ;
  LAYER metal2 ;
  RECT 0.000 901.940 1.120 905.180 ;
  LAYER metal1 ;
  RECT 0.000 901.940 1.120 905.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 894.100 1.120 897.340 ;
  LAYER metal3 ;
  RECT 0.000 894.100 1.120 897.340 ;
  LAYER metal2 ;
  RECT 0.000 894.100 1.120 897.340 ;
  LAYER metal1 ;
  RECT 0.000 894.100 1.120 897.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 886.260 1.120 889.500 ;
  LAYER metal3 ;
  RECT 0.000 886.260 1.120 889.500 ;
  LAYER metal2 ;
  RECT 0.000 886.260 1.120 889.500 ;
  LAYER metal1 ;
  RECT 0.000 886.260 1.120 889.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 878.420 1.120 881.660 ;
  LAYER metal3 ;
  RECT 0.000 878.420 1.120 881.660 ;
  LAYER metal2 ;
  RECT 0.000 878.420 1.120 881.660 ;
  LAYER metal1 ;
  RECT 0.000 878.420 1.120 881.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 870.580 1.120 873.820 ;
  LAYER metal3 ;
  RECT 0.000 870.580 1.120 873.820 ;
  LAYER metal2 ;
  RECT 0.000 870.580 1.120 873.820 ;
  LAYER metal1 ;
  RECT 0.000 870.580 1.120 873.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 831.380 1.120 834.620 ;
  LAYER metal3 ;
  RECT 0.000 831.380 1.120 834.620 ;
  LAYER metal2 ;
  RECT 0.000 831.380 1.120 834.620 ;
  LAYER metal1 ;
  RECT 0.000 831.380 1.120 834.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 823.540 1.120 826.780 ;
  LAYER metal3 ;
  RECT 0.000 823.540 1.120 826.780 ;
  LAYER metal2 ;
  RECT 0.000 823.540 1.120 826.780 ;
  LAYER metal1 ;
  RECT 0.000 823.540 1.120 826.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 815.700 1.120 818.940 ;
  LAYER metal3 ;
  RECT 0.000 815.700 1.120 818.940 ;
  LAYER metal2 ;
  RECT 0.000 815.700 1.120 818.940 ;
  LAYER metal1 ;
  RECT 0.000 815.700 1.120 818.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 807.860 1.120 811.100 ;
  LAYER metal3 ;
  RECT 0.000 807.860 1.120 811.100 ;
  LAYER metal2 ;
  RECT 0.000 807.860 1.120 811.100 ;
  LAYER metal1 ;
  RECT 0.000 807.860 1.120 811.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 800.020 1.120 803.260 ;
  LAYER metal3 ;
  RECT 0.000 800.020 1.120 803.260 ;
  LAYER metal2 ;
  RECT 0.000 800.020 1.120 803.260 ;
  LAYER metal1 ;
  RECT 0.000 800.020 1.120 803.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 792.180 1.120 795.420 ;
  LAYER metal3 ;
  RECT 0.000 792.180 1.120 795.420 ;
  LAYER metal2 ;
  RECT 0.000 792.180 1.120 795.420 ;
  LAYER metal1 ;
  RECT 0.000 792.180 1.120 795.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 752.980 1.120 756.220 ;
  LAYER metal3 ;
  RECT 0.000 752.980 1.120 756.220 ;
  LAYER metal2 ;
  RECT 0.000 752.980 1.120 756.220 ;
  LAYER metal1 ;
  RECT 0.000 752.980 1.120 756.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 745.140 1.120 748.380 ;
  LAYER metal3 ;
  RECT 0.000 745.140 1.120 748.380 ;
  LAYER metal2 ;
  RECT 0.000 745.140 1.120 748.380 ;
  LAYER metal1 ;
  RECT 0.000 745.140 1.120 748.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 737.300 1.120 740.540 ;
  LAYER metal3 ;
  RECT 0.000 737.300 1.120 740.540 ;
  LAYER metal2 ;
  RECT 0.000 737.300 1.120 740.540 ;
  LAYER metal1 ;
  RECT 0.000 737.300 1.120 740.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 729.460 1.120 732.700 ;
  LAYER metal3 ;
  RECT 0.000 729.460 1.120 732.700 ;
  LAYER metal2 ;
  RECT 0.000 729.460 1.120 732.700 ;
  LAYER metal1 ;
  RECT 0.000 729.460 1.120 732.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 721.620 1.120 724.860 ;
  LAYER metal3 ;
  RECT 0.000 721.620 1.120 724.860 ;
  LAYER metal2 ;
  RECT 0.000 721.620 1.120 724.860 ;
  LAYER metal1 ;
  RECT 0.000 721.620 1.120 724.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 713.780 1.120 717.020 ;
  LAYER metal3 ;
  RECT 0.000 713.780 1.120 717.020 ;
  LAYER metal2 ;
  RECT 0.000 713.780 1.120 717.020 ;
  LAYER metal1 ;
  RECT 0.000 713.780 1.120 717.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 674.580 1.120 677.820 ;
  LAYER metal3 ;
  RECT 0.000 674.580 1.120 677.820 ;
  LAYER metal2 ;
  RECT 0.000 674.580 1.120 677.820 ;
  LAYER metal1 ;
  RECT 0.000 674.580 1.120 677.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 666.740 1.120 669.980 ;
  LAYER metal3 ;
  RECT 0.000 666.740 1.120 669.980 ;
  LAYER metal2 ;
  RECT 0.000 666.740 1.120 669.980 ;
  LAYER metal1 ;
  RECT 0.000 666.740 1.120 669.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 658.900 1.120 662.140 ;
  LAYER metal3 ;
  RECT 0.000 658.900 1.120 662.140 ;
  LAYER metal2 ;
  RECT 0.000 658.900 1.120 662.140 ;
  LAYER metal1 ;
  RECT 0.000 658.900 1.120 662.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 651.060 1.120 654.300 ;
  LAYER metal3 ;
  RECT 0.000 651.060 1.120 654.300 ;
  LAYER metal2 ;
  RECT 0.000 651.060 1.120 654.300 ;
  LAYER metal1 ;
  RECT 0.000 651.060 1.120 654.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 643.220 1.120 646.460 ;
  LAYER metal3 ;
  RECT 0.000 643.220 1.120 646.460 ;
  LAYER metal2 ;
  RECT 0.000 643.220 1.120 646.460 ;
  LAYER metal1 ;
  RECT 0.000 643.220 1.120 646.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 635.380 1.120 638.620 ;
  LAYER metal3 ;
  RECT 0.000 635.380 1.120 638.620 ;
  LAYER metal2 ;
  RECT 0.000 635.380 1.120 638.620 ;
  LAYER metal1 ;
  RECT 0.000 635.380 1.120 638.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 596.180 1.120 599.420 ;
  LAYER metal3 ;
  RECT 0.000 596.180 1.120 599.420 ;
  LAYER metal2 ;
  RECT 0.000 596.180 1.120 599.420 ;
  LAYER metal1 ;
  RECT 0.000 596.180 1.120 599.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 588.340 1.120 591.580 ;
  LAYER metal3 ;
  RECT 0.000 588.340 1.120 591.580 ;
  LAYER metal2 ;
  RECT 0.000 588.340 1.120 591.580 ;
  LAYER metal1 ;
  RECT 0.000 588.340 1.120 591.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 580.500 1.120 583.740 ;
  LAYER metal3 ;
  RECT 0.000 580.500 1.120 583.740 ;
  LAYER metal2 ;
  RECT 0.000 580.500 1.120 583.740 ;
  LAYER metal1 ;
  RECT 0.000 580.500 1.120 583.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 572.660 1.120 575.900 ;
  LAYER metal3 ;
  RECT 0.000 572.660 1.120 575.900 ;
  LAYER metal2 ;
  RECT 0.000 572.660 1.120 575.900 ;
  LAYER metal1 ;
  RECT 0.000 572.660 1.120 575.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 564.820 1.120 568.060 ;
  LAYER metal3 ;
  RECT 0.000 564.820 1.120 568.060 ;
  LAYER metal2 ;
  RECT 0.000 564.820 1.120 568.060 ;
  LAYER metal1 ;
  RECT 0.000 564.820 1.120 568.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 556.980 1.120 560.220 ;
  LAYER metal3 ;
  RECT 0.000 556.980 1.120 560.220 ;
  LAYER metal2 ;
  RECT 0.000 556.980 1.120 560.220 ;
  LAYER metal1 ;
  RECT 0.000 556.980 1.120 560.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER metal3 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER metal2 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER metal1 ;
  RECT 0.000 517.780 1.120 521.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER metal3 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER metal2 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER metal1 ;
  RECT 0.000 509.940 1.120 513.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER metal3 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER metal2 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER metal1 ;
  RECT 0.000 502.100 1.120 505.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER metal3 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER metal2 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER metal1 ;
  RECT 0.000 494.260 1.120 497.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER metal3 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER metal2 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER metal1 ;
  RECT 0.000 486.420 1.120 489.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER metal3 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER metal2 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER metal1 ;
  RECT 0.000 478.580 1.120 481.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER metal3 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER metal2 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER metal1 ;
  RECT 0.000 439.380 1.120 442.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER metal3 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER metal2 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER metal1 ;
  RECT 0.000 431.540 1.120 434.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER metal3 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER metal2 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER metal1 ;
  RECT 0.000 423.700 1.120 426.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER metal3 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER metal2 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER metal1 ;
  RECT 0.000 415.860 1.120 419.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER metal3 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER metal2 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER metal1 ;
  RECT 0.000 408.020 1.120 411.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER metal3 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER metal2 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER metal1 ;
  RECT 0.000 400.180 1.120 403.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER metal3 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER metal2 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER metal1 ;
  RECT 0.000 360.980 1.120 364.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER metal3 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER metal2 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER metal1 ;
  RECT 0.000 353.140 1.120 356.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER metal3 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER metal2 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER metal1 ;
  RECT 0.000 345.300 1.120 348.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER metal3 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER metal2 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER metal1 ;
  RECT 0.000 337.460 1.120 340.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER metal3 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER metal2 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER metal1 ;
  RECT 0.000 329.620 1.120 332.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER metal3 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER metal2 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER metal1 ;
  RECT 0.000 321.780 1.120 325.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal3 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal2 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal1 ;
  RECT 0.000 282.580 1.120 285.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal3 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal2 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal1 ;
  RECT 0.000 274.740 1.120 277.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal3 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal2 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal1 ;
  RECT 0.000 266.900 1.120 270.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal3 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal2 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal1 ;
  RECT 0.000 259.060 1.120 262.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal3 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal2 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal1 ;
  RECT 0.000 251.220 1.120 254.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal3 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal2 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal1 ;
  RECT 0.000 243.380 1.120 246.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1874.040 1390.480 1877.580 1391.600 ;
  LAYER metal3 ;
  RECT 1874.040 1390.480 1877.580 1391.600 ;
  LAYER metal2 ;
  RECT 1874.040 1390.480 1877.580 1391.600 ;
  LAYER metal1 ;
  RECT 1874.040 1390.480 1877.580 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1865.360 1390.480 1868.900 1391.600 ;
  LAYER metal3 ;
  RECT 1865.360 1390.480 1868.900 1391.600 ;
  LAYER metal2 ;
  RECT 1865.360 1390.480 1868.900 1391.600 ;
  LAYER metal1 ;
  RECT 1865.360 1390.480 1868.900 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1856.680 1390.480 1860.220 1391.600 ;
  LAYER metal3 ;
  RECT 1856.680 1390.480 1860.220 1391.600 ;
  LAYER metal2 ;
  RECT 1856.680 1390.480 1860.220 1391.600 ;
  LAYER metal1 ;
  RECT 1856.680 1390.480 1860.220 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1848.000 1390.480 1851.540 1391.600 ;
  LAYER metal3 ;
  RECT 1848.000 1390.480 1851.540 1391.600 ;
  LAYER metal2 ;
  RECT 1848.000 1390.480 1851.540 1391.600 ;
  LAYER metal1 ;
  RECT 1848.000 1390.480 1851.540 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1839.320 1390.480 1842.860 1391.600 ;
  LAYER metal3 ;
  RECT 1839.320 1390.480 1842.860 1391.600 ;
  LAYER metal2 ;
  RECT 1839.320 1390.480 1842.860 1391.600 ;
  LAYER metal1 ;
  RECT 1839.320 1390.480 1842.860 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1830.640 1390.480 1834.180 1391.600 ;
  LAYER metal3 ;
  RECT 1830.640 1390.480 1834.180 1391.600 ;
  LAYER metal2 ;
  RECT 1830.640 1390.480 1834.180 1391.600 ;
  LAYER metal1 ;
  RECT 1830.640 1390.480 1834.180 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1787.240 1390.480 1790.780 1391.600 ;
  LAYER metal3 ;
  RECT 1787.240 1390.480 1790.780 1391.600 ;
  LAYER metal2 ;
  RECT 1787.240 1390.480 1790.780 1391.600 ;
  LAYER metal1 ;
  RECT 1787.240 1390.480 1790.780 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1778.560 1390.480 1782.100 1391.600 ;
  LAYER metal3 ;
  RECT 1778.560 1390.480 1782.100 1391.600 ;
  LAYER metal2 ;
  RECT 1778.560 1390.480 1782.100 1391.600 ;
  LAYER metal1 ;
  RECT 1778.560 1390.480 1782.100 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1769.880 1390.480 1773.420 1391.600 ;
  LAYER metal3 ;
  RECT 1769.880 1390.480 1773.420 1391.600 ;
  LAYER metal2 ;
  RECT 1769.880 1390.480 1773.420 1391.600 ;
  LAYER metal1 ;
  RECT 1769.880 1390.480 1773.420 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1761.200 1390.480 1764.740 1391.600 ;
  LAYER metal3 ;
  RECT 1761.200 1390.480 1764.740 1391.600 ;
  LAYER metal2 ;
  RECT 1761.200 1390.480 1764.740 1391.600 ;
  LAYER metal1 ;
  RECT 1761.200 1390.480 1764.740 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1752.520 1390.480 1756.060 1391.600 ;
  LAYER metal3 ;
  RECT 1752.520 1390.480 1756.060 1391.600 ;
  LAYER metal2 ;
  RECT 1752.520 1390.480 1756.060 1391.600 ;
  LAYER metal1 ;
  RECT 1752.520 1390.480 1756.060 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1743.840 1390.480 1747.380 1391.600 ;
  LAYER metal3 ;
  RECT 1743.840 1390.480 1747.380 1391.600 ;
  LAYER metal2 ;
  RECT 1743.840 1390.480 1747.380 1391.600 ;
  LAYER metal1 ;
  RECT 1743.840 1390.480 1747.380 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1700.440 1390.480 1703.980 1391.600 ;
  LAYER metal3 ;
  RECT 1700.440 1390.480 1703.980 1391.600 ;
  LAYER metal2 ;
  RECT 1700.440 1390.480 1703.980 1391.600 ;
  LAYER metal1 ;
  RECT 1700.440 1390.480 1703.980 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1691.760 1390.480 1695.300 1391.600 ;
  LAYER metal3 ;
  RECT 1691.760 1390.480 1695.300 1391.600 ;
  LAYER metal2 ;
  RECT 1691.760 1390.480 1695.300 1391.600 ;
  LAYER metal1 ;
  RECT 1691.760 1390.480 1695.300 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1683.080 1390.480 1686.620 1391.600 ;
  LAYER metal3 ;
  RECT 1683.080 1390.480 1686.620 1391.600 ;
  LAYER metal2 ;
  RECT 1683.080 1390.480 1686.620 1391.600 ;
  LAYER metal1 ;
  RECT 1683.080 1390.480 1686.620 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1674.400 1390.480 1677.940 1391.600 ;
  LAYER metal3 ;
  RECT 1674.400 1390.480 1677.940 1391.600 ;
  LAYER metal2 ;
  RECT 1674.400 1390.480 1677.940 1391.600 ;
  LAYER metal1 ;
  RECT 1674.400 1390.480 1677.940 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1665.720 1390.480 1669.260 1391.600 ;
  LAYER metal3 ;
  RECT 1665.720 1390.480 1669.260 1391.600 ;
  LAYER metal2 ;
  RECT 1665.720 1390.480 1669.260 1391.600 ;
  LAYER metal1 ;
  RECT 1665.720 1390.480 1669.260 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1657.040 1390.480 1660.580 1391.600 ;
  LAYER metal3 ;
  RECT 1657.040 1390.480 1660.580 1391.600 ;
  LAYER metal2 ;
  RECT 1657.040 1390.480 1660.580 1391.600 ;
  LAYER metal1 ;
  RECT 1657.040 1390.480 1660.580 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1613.640 1390.480 1617.180 1391.600 ;
  LAYER metal3 ;
  RECT 1613.640 1390.480 1617.180 1391.600 ;
  LAYER metal2 ;
  RECT 1613.640 1390.480 1617.180 1391.600 ;
  LAYER metal1 ;
  RECT 1613.640 1390.480 1617.180 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1604.960 1390.480 1608.500 1391.600 ;
  LAYER metal3 ;
  RECT 1604.960 1390.480 1608.500 1391.600 ;
  LAYER metal2 ;
  RECT 1604.960 1390.480 1608.500 1391.600 ;
  LAYER metal1 ;
  RECT 1604.960 1390.480 1608.500 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1596.280 1390.480 1599.820 1391.600 ;
  LAYER metal3 ;
  RECT 1596.280 1390.480 1599.820 1391.600 ;
  LAYER metal2 ;
  RECT 1596.280 1390.480 1599.820 1391.600 ;
  LAYER metal1 ;
  RECT 1596.280 1390.480 1599.820 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1587.600 1390.480 1591.140 1391.600 ;
  LAYER metal3 ;
  RECT 1587.600 1390.480 1591.140 1391.600 ;
  LAYER metal2 ;
  RECT 1587.600 1390.480 1591.140 1391.600 ;
  LAYER metal1 ;
  RECT 1587.600 1390.480 1591.140 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1578.920 1390.480 1582.460 1391.600 ;
  LAYER metal3 ;
  RECT 1578.920 1390.480 1582.460 1391.600 ;
  LAYER metal2 ;
  RECT 1578.920 1390.480 1582.460 1391.600 ;
  LAYER metal1 ;
  RECT 1578.920 1390.480 1582.460 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1570.240 1390.480 1573.780 1391.600 ;
  LAYER metal3 ;
  RECT 1570.240 1390.480 1573.780 1391.600 ;
  LAYER metal2 ;
  RECT 1570.240 1390.480 1573.780 1391.600 ;
  LAYER metal1 ;
  RECT 1570.240 1390.480 1573.780 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1526.840 1390.480 1530.380 1391.600 ;
  LAYER metal3 ;
  RECT 1526.840 1390.480 1530.380 1391.600 ;
  LAYER metal2 ;
  RECT 1526.840 1390.480 1530.380 1391.600 ;
  LAYER metal1 ;
  RECT 1526.840 1390.480 1530.380 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1518.160 1390.480 1521.700 1391.600 ;
  LAYER metal3 ;
  RECT 1518.160 1390.480 1521.700 1391.600 ;
  LAYER metal2 ;
  RECT 1518.160 1390.480 1521.700 1391.600 ;
  LAYER metal1 ;
  RECT 1518.160 1390.480 1521.700 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1509.480 1390.480 1513.020 1391.600 ;
  LAYER metal3 ;
  RECT 1509.480 1390.480 1513.020 1391.600 ;
  LAYER metal2 ;
  RECT 1509.480 1390.480 1513.020 1391.600 ;
  LAYER metal1 ;
  RECT 1509.480 1390.480 1513.020 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1500.800 1390.480 1504.340 1391.600 ;
  LAYER metal3 ;
  RECT 1500.800 1390.480 1504.340 1391.600 ;
  LAYER metal2 ;
  RECT 1500.800 1390.480 1504.340 1391.600 ;
  LAYER metal1 ;
  RECT 1500.800 1390.480 1504.340 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1492.120 1390.480 1495.660 1391.600 ;
  LAYER metal3 ;
  RECT 1492.120 1390.480 1495.660 1391.600 ;
  LAYER metal2 ;
  RECT 1492.120 1390.480 1495.660 1391.600 ;
  LAYER metal1 ;
  RECT 1492.120 1390.480 1495.660 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1483.440 1390.480 1486.980 1391.600 ;
  LAYER metal3 ;
  RECT 1483.440 1390.480 1486.980 1391.600 ;
  LAYER metal2 ;
  RECT 1483.440 1390.480 1486.980 1391.600 ;
  LAYER metal1 ;
  RECT 1483.440 1390.480 1486.980 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1440.040 1390.480 1443.580 1391.600 ;
  LAYER metal3 ;
  RECT 1440.040 1390.480 1443.580 1391.600 ;
  LAYER metal2 ;
  RECT 1440.040 1390.480 1443.580 1391.600 ;
  LAYER metal1 ;
  RECT 1440.040 1390.480 1443.580 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1431.360 1390.480 1434.900 1391.600 ;
  LAYER metal3 ;
  RECT 1431.360 1390.480 1434.900 1391.600 ;
  LAYER metal2 ;
  RECT 1431.360 1390.480 1434.900 1391.600 ;
  LAYER metal1 ;
  RECT 1431.360 1390.480 1434.900 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1422.680 1390.480 1426.220 1391.600 ;
  LAYER metal3 ;
  RECT 1422.680 1390.480 1426.220 1391.600 ;
  LAYER metal2 ;
  RECT 1422.680 1390.480 1426.220 1391.600 ;
  LAYER metal1 ;
  RECT 1422.680 1390.480 1426.220 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1414.000 1390.480 1417.540 1391.600 ;
  LAYER metal3 ;
  RECT 1414.000 1390.480 1417.540 1391.600 ;
  LAYER metal2 ;
  RECT 1414.000 1390.480 1417.540 1391.600 ;
  LAYER metal1 ;
  RECT 1414.000 1390.480 1417.540 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1405.320 1390.480 1408.860 1391.600 ;
  LAYER metal3 ;
  RECT 1405.320 1390.480 1408.860 1391.600 ;
  LAYER metal2 ;
  RECT 1405.320 1390.480 1408.860 1391.600 ;
  LAYER metal1 ;
  RECT 1405.320 1390.480 1408.860 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1396.640 1390.480 1400.180 1391.600 ;
  LAYER metal3 ;
  RECT 1396.640 1390.480 1400.180 1391.600 ;
  LAYER metal2 ;
  RECT 1396.640 1390.480 1400.180 1391.600 ;
  LAYER metal1 ;
  RECT 1396.640 1390.480 1400.180 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1353.240 1390.480 1356.780 1391.600 ;
  LAYER metal3 ;
  RECT 1353.240 1390.480 1356.780 1391.600 ;
  LAYER metal2 ;
  RECT 1353.240 1390.480 1356.780 1391.600 ;
  LAYER metal1 ;
  RECT 1353.240 1390.480 1356.780 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1344.560 1390.480 1348.100 1391.600 ;
  LAYER metal3 ;
  RECT 1344.560 1390.480 1348.100 1391.600 ;
  LAYER metal2 ;
  RECT 1344.560 1390.480 1348.100 1391.600 ;
  LAYER metal1 ;
  RECT 1344.560 1390.480 1348.100 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1335.880 1390.480 1339.420 1391.600 ;
  LAYER metal3 ;
  RECT 1335.880 1390.480 1339.420 1391.600 ;
  LAYER metal2 ;
  RECT 1335.880 1390.480 1339.420 1391.600 ;
  LAYER metal1 ;
  RECT 1335.880 1390.480 1339.420 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1327.200 1390.480 1330.740 1391.600 ;
  LAYER metal3 ;
  RECT 1327.200 1390.480 1330.740 1391.600 ;
  LAYER metal2 ;
  RECT 1327.200 1390.480 1330.740 1391.600 ;
  LAYER metal1 ;
  RECT 1327.200 1390.480 1330.740 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1318.520 1390.480 1322.060 1391.600 ;
  LAYER metal3 ;
  RECT 1318.520 1390.480 1322.060 1391.600 ;
  LAYER metal2 ;
  RECT 1318.520 1390.480 1322.060 1391.600 ;
  LAYER metal1 ;
  RECT 1318.520 1390.480 1322.060 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1309.840 1390.480 1313.380 1391.600 ;
  LAYER metal3 ;
  RECT 1309.840 1390.480 1313.380 1391.600 ;
  LAYER metal2 ;
  RECT 1309.840 1390.480 1313.380 1391.600 ;
  LAYER metal1 ;
  RECT 1309.840 1390.480 1313.380 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1266.440 1390.480 1269.980 1391.600 ;
  LAYER metal3 ;
  RECT 1266.440 1390.480 1269.980 1391.600 ;
  LAYER metal2 ;
  RECT 1266.440 1390.480 1269.980 1391.600 ;
  LAYER metal1 ;
  RECT 1266.440 1390.480 1269.980 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1257.760 1390.480 1261.300 1391.600 ;
  LAYER metal3 ;
  RECT 1257.760 1390.480 1261.300 1391.600 ;
  LAYER metal2 ;
  RECT 1257.760 1390.480 1261.300 1391.600 ;
  LAYER metal1 ;
  RECT 1257.760 1390.480 1261.300 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1249.080 1390.480 1252.620 1391.600 ;
  LAYER metal3 ;
  RECT 1249.080 1390.480 1252.620 1391.600 ;
  LAYER metal2 ;
  RECT 1249.080 1390.480 1252.620 1391.600 ;
  LAYER metal1 ;
  RECT 1249.080 1390.480 1252.620 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1240.400 1390.480 1243.940 1391.600 ;
  LAYER metal3 ;
  RECT 1240.400 1390.480 1243.940 1391.600 ;
  LAYER metal2 ;
  RECT 1240.400 1390.480 1243.940 1391.600 ;
  LAYER metal1 ;
  RECT 1240.400 1390.480 1243.940 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1231.720 1390.480 1235.260 1391.600 ;
  LAYER metal3 ;
  RECT 1231.720 1390.480 1235.260 1391.600 ;
  LAYER metal2 ;
  RECT 1231.720 1390.480 1235.260 1391.600 ;
  LAYER metal1 ;
  RECT 1231.720 1390.480 1235.260 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1223.040 1390.480 1226.580 1391.600 ;
  LAYER metal3 ;
  RECT 1223.040 1390.480 1226.580 1391.600 ;
  LAYER metal2 ;
  RECT 1223.040 1390.480 1226.580 1391.600 ;
  LAYER metal1 ;
  RECT 1223.040 1390.480 1226.580 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1179.640 1390.480 1183.180 1391.600 ;
  LAYER metal3 ;
  RECT 1179.640 1390.480 1183.180 1391.600 ;
  LAYER metal2 ;
  RECT 1179.640 1390.480 1183.180 1391.600 ;
  LAYER metal1 ;
  RECT 1179.640 1390.480 1183.180 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1170.960 1390.480 1174.500 1391.600 ;
  LAYER metal3 ;
  RECT 1170.960 1390.480 1174.500 1391.600 ;
  LAYER metal2 ;
  RECT 1170.960 1390.480 1174.500 1391.600 ;
  LAYER metal1 ;
  RECT 1170.960 1390.480 1174.500 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1162.280 1390.480 1165.820 1391.600 ;
  LAYER metal3 ;
  RECT 1162.280 1390.480 1165.820 1391.600 ;
  LAYER metal2 ;
  RECT 1162.280 1390.480 1165.820 1391.600 ;
  LAYER metal1 ;
  RECT 1162.280 1390.480 1165.820 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1153.600 1390.480 1157.140 1391.600 ;
  LAYER metal3 ;
  RECT 1153.600 1390.480 1157.140 1391.600 ;
  LAYER metal2 ;
  RECT 1153.600 1390.480 1157.140 1391.600 ;
  LAYER metal1 ;
  RECT 1153.600 1390.480 1157.140 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1144.920 1390.480 1148.460 1391.600 ;
  LAYER metal3 ;
  RECT 1144.920 1390.480 1148.460 1391.600 ;
  LAYER metal2 ;
  RECT 1144.920 1390.480 1148.460 1391.600 ;
  LAYER metal1 ;
  RECT 1144.920 1390.480 1148.460 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1136.240 1390.480 1139.780 1391.600 ;
  LAYER metal3 ;
  RECT 1136.240 1390.480 1139.780 1391.600 ;
  LAYER metal2 ;
  RECT 1136.240 1390.480 1139.780 1391.600 ;
  LAYER metal1 ;
  RECT 1136.240 1390.480 1139.780 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1092.840 1390.480 1096.380 1391.600 ;
  LAYER metal3 ;
  RECT 1092.840 1390.480 1096.380 1391.600 ;
  LAYER metal2 ;
  RECT 1092.840 1390.480 1096.380 1391.600 ;
  LAYER metal1 ;
  RECT 1092.840 1390.480 1096.380 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1084.160 1390.480 1087.700 1391.600 ;
  LAYER metal3 ;
  RECT 1084.160 1390.480 1087.700 1391.600 ;
  LAYER metal2 ;
  RECT 1084.160 1390.480 1087.700 1391.600 ;
  LAYER metal1 ;
  RECT 1084.160 1390.480 1087.700 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1075.480 1390.480 1079.020 1391.600 ;
  LAYER metal3 ;
  RECT 1075.480 1390.480 1079.020 1391.600 ;
  LAYER metal2 ;
  RECT 1075.480 1390.480 1079.020 1391.600 ;
  LAYER metal1 ;
  RECT 1075.480 1390.480 1079.020 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1066.800 1390.480 1070.340 1391.600 ;
  LAYER metal3 ;
  RECT 1066.800 1390.480 1070.340 1391.600 ;
  LAYER metal2 ;
  RECT 1066.800 1390.480 1070.340 1391.600 ;
  LAYER metal1 ;
  RECT 1066.800 1390.480 1070.340 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1058.120 1390.480 1061.660 1391.600 ;
  LAYER metal3 ;
  RECT 1058.120 1390.480 1061.660 1391.600 ;
  LAYER metal2 ;
  RECT 1058.120 1390.480 1061.660 1391.600 ;
  LAYER metal1 ;
  RECT 1058.120 1390.480 1061.660 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1049.440 1390.480 1052.980 1391.600 ;
  LAYER metal3 ;
  RECT 1049.440 1390.480 1052.980 1391.600 ;
  LAYER metal2 ;
  RECT 1049.440 1390.480 1052.980 1391.600 ;
  LAYER metal1 ;
  RECT 1049.440 1390.480 1052.980 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1006.040 1390.480 1009.580 1391.600 ;
  LAYER metal3 ;
  RECT 1006.040 1390.480 1009.580 1391.600 ;
  LAYER metal2 ;
  RECT 1006.040 1390.480 1009.580 1391.600 ;
  LAYER metal1 ;
  RECT 1006.040 1390.480 1009.580 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 997.360 1390.480 1000.900 1391.600 ;
  LAYER metal3 ;
  RECT 997.360 1390.480 1000.900 1391.600 ;
  LAYER metal2 ;
  RECT 997.360 1390.480 1000.900 1391.600 ;
  LAYER metal1 ;
  RECT 997.360 1390.480 1000.900 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 988.680 1390.480 992.220 1391.600 ;
  LAYER metal3 ;
  RECT 988.680 1390.480 992.220 1391.600 ;
  LAYER metal2 ;
  RECT 988.680 1390.480 992.220 1391.600 ;
  LAYER metal1 ;
  RECT 988.680 1390.480 992.220 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 980.000 1390.480 983.540 1391.600 ;
  LAYER metal3 ;
  RECT 980.000 1390.480 983.540 1391.600 ;
  LAYER metal2 ;
  RECT 980.000 1390.480 983.540 1391.600 ;
  LAYER metal1 ;
  RECT 980.000 1390.480 983.540 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 971.320 1390.480 974.860 1391.600 ;
  LAYER metal3 ;
  RECT 971.320 1390.480 974.860 1391.600 ;
  LAYER metal2 ;
  RECT 971.320 1390.480 974.860 1391.600 ;
  LAYER metal1 ;
  RECT 971.320 1390.480 974.860 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 962.640 1390.480 966.180 1391.600 ;
  LAYER metal3 ;
  RECT 962.640 1390.480 966.180 1391.600 ;
  LAYER metal2 ;
  RECT 962.640 1390.480 966.180 1391.600 ;
  LAYER metal1 ;
  RECT 962.640 1390.480 966.180 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 919.240 1390.480 922.780 1391.600 ;
  LAYER metal3 ;
  RECT 919.240 1390.480 922.780 1391.600 ;
  LAYER metal2 ;
  RECT 919.240 1390.480 922.780 1391.600 ;
  LAYER metal1 ;
  RECT 919.240 1390.480 922.780 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 910.560 1390.480 914.100 1391.600 ;
  LAYER metal3 ;
  RECT 910.560 1390.480 914.100 1391.600 ;
  LAYER metal2 ;
  RECT 910.560 1390.480 914.100 1391.600 ;
  LAYER metal1 ;
  RECT 910.560 1390.480 914.100 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 901.880 1390.480 905.420 1391.600 ;
  LAYER metal3 ;
  RECT 901.880 1390.480 905.420 1391.600 ;
  LAYER metal2 ;
  RECT 901.880 1390.480 905.420 1391.600 ;
  LAYER metal1 ;
  RECT 901.880 1390.480 905.420 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 893.200 1390.480 896.740 1391.600 ;
  LAYER metal3 ;
  RECT 893.200 1390.480 896.740 1391.600 ;
  LAYER metal2 ;
  RECT 893.200 1390.480 896.740 1391.600 ;
  LAYER metal1 ;
  RECT 893.200 1390.480 896.740 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 884.520 1390.480 888.060 1391.600 ;
  LAYER metal3 ;
  RECT 884.520 1390.480 888.060 1391.600 ;
  LAYER metal2 ;
  RECT 884.520 1390.480 888.060 1391.600 ;
  LAYER metal1 ;
  RECT 884.520 1390.480 888.060 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 875.840 1390.480 879.380 1391.600 ;
  LAYER metal3 ;
  RECT 875.840 1390.480 879.380 1391.600 ;
  LAYER metal2 ;
  RECT 875.840 1390.480 879.380 1391.600 ;
  LAYER metal1 ;
  RECT 875.840 1390.480 879.380 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 832.440 1390.480 835.980 1391.600 ;
  LAYER metal3 ;
  RECT 832.440 1390.480 835.980 1391.600 ;
  LAYER metal2 ;
  RECT 832.440 1390.480 835.980 1391.600 ;
  LAYER metal1 ;
  RECT 832.440 1390.480 835.980 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 823.760 1390.480 827.300 1391.600 ;
  LAYER metal3 ;
  RECT 823.760 1390.480 827.300 1391.600 ;
  LAYER metal2 ;
  RECT 823.760 1390.480 827.300 1391.600 ;
  LAYER metal1 ;
  RECT 823.760 1390.480 827.300 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 815.080 1390.480 818.620 1391.600 ;
  LAYER metal3 ;
  RECT 815.080 1390.480 818.620 1391.600 ;
  LAYER metal2 ;
  RECT 815.080 1390.480 818.620 1391.600 ;
  LAYER metal1 ;
  RECT 815.080 1390.480 818.620 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 806.400 1390.480 809.940 1391.600 ;
  LAYER metal3 ;
  RECT 806.400 1390.480 809.940 1391.600 ;
  LAYER metal2 ;
  RECT 806.400 1390.480 809.940 1391.600 ;
  LAYER metal1 ;
  RECT 806.400 1390.480 809.940 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 797.720 1390.480 801.260 1391.600 ;
  LAYER metal3 ;
  RECT 797.720 1390.480 801.260 1391.600 ;
  LAYER metal2 ;
  RECT 797.720 1390.480 801.260 1391.600 ;
  LAYER metal1 ;
  RECT 797.720 1390.480 801.260 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 789.040 1390.480 792.580 1391.600 ;
  LAYER metal3 ;
  RECT 789.040 1390.480 792.580 1391.600 ;
  LAYER metal2 ;
  RECT 789.040 1390.480 792.580 1391.600 ;
  LAYER metal1 ;
  RECT 789.040 1390.480 792.580 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 745.640 1390.480 749.180 1391.600 ;
  LAYER metal3 ;
  RECT 745.640 1390.480 749.180 1391.600 ;
  LAYER metal2 ;
  RECT 745.640 1390.480 749.180 1391.600 ;
  LAYER metal1 ;
  RECT 745.640 1390.480 749.180 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 736.960 1390.480 740.500 1391.600 ;
  LAYER metal3 ;
  RECT 736.960 1390.480 740.500 1391.600 ;
  LAYER metal2 ;
  RECT 736.960 1390.480 740.500 1391.600 ;
  LAYER metal1 ;
  RECT 736.960 1390.480 740.500 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 728.280 1390.480 731.820 1391.600 ;
  LAYER metal3 ;
  RECT 728.280 1390.480 731.820 1391.600 ;
  LAYER metal2 ;
  RECT 728.280 1390.480 731.820 1391.600 ;
  LAYER metal1 ;
  RECT 728.280 1390.480 731.820 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 719.600 1390.480 723.140 1391.600 ;
  LAYER metal3 ;
  RECT 719.600 1390.480 723.140 1391.600 ;
  LAYER metal2 ;
  RECT 719.600 1390.480 723.140 1391.600 ;
  LAYER metal1 ;
  RECT 719.600 1390.480 723.140 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 710.920 1390.480 714.460 1391.600 ;
  LAYER metal3 ;
  RECT 710.920 1390.480 714.460 1391.600 ;
  LAYER metal2 ;
  RECT 710.920 1390.480 714.460 1391.600 ;
  LAYER metal1 ;
  RECT 710.920 1390.480 714.460 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 702.240 1390.480 705.780 1391.600 ;
  LAYER metal3 ;
  RECT 702.240 1390.480 705.780 1391.600 ;
  LAYER metal2 ;
  RECT 702.240 1390.480 705.780 1391.600 ;
  LAYER metal1 ;
  RECT 702.240 1390.480 705.780 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 658.840 1390.480 662.380 1391.600 ;
  LAYER metal3 ;
  RECT 658.840 1390.480 662.380 1391.600 ;
  LAYER metal2 ;
  RECT 658.840 1390.480 662.380 1391.600 ;
  LAYER metal1 ;
  RECT 658.840 1390.480 662.380 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 650.160 1390.480 653.700 1391.600 ;
  LAYER metal3 ;
  RECT 650.160 1390.480 653.700 1391.600 ;
  LAYER metal2 ;
  RECT 650.160 1390.480 653.700 1391.600 ;
  LAYER metal1 ;
  RECT 650.160 1390.480 653.700 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 641.480 1390.480 645.020 1391.600 ;
  LAYER metal3 ;
  RECT 641.480 1390.480 645.020 1391.600 ;
  LAYER metal2 ;
  RECT 641.480 1390.480 645.020 1391.600 ;
  LAYER metal1 ;
  RECT 641.480 1390.480 645.020 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 632.800 1390.480 636.340 1391.600 ;
  LAYER metal3 ;
  RECT 632.800 1390.480 636.340 1391.600 ;
  LAYER metal2 ;
  RECT 632.800 1390.480 636.340 1391.600 ;
  LAYER metal1 ;
  RECT 632.800 1390.480 636.340 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 624.120 1390.480 627.660 1391.600 ;
  LAYER metal3 ;
  RECT 624.120 1390.480 627.660 1391.600 ;
  LAYER metal2 ;
  RECT 624.120 1390.480 627.660 1391.600 ;
  LAYER metal1 ;
  RECT 624.120 1390.480 627.660 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 615.440 1390.480 618.980 1391.600 ;
  LAYER metal3 ;
  RECT 615.440 1390.480 618.980 1391.600 ;
  LAYER metal2 ;
  RECT 615.440 1390.480 618.980 1391.600 ;
  LAYER metal1 ;
  RECT 615.440 1390.480 618.980 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 572.040 1390.480 575.580 1391.600 ;
  LAYER metal3 ;
  RECT 572.040 1390.480 575.580 1391.600 ;
  LAYER metal2 ;
  RECT 572.040 1390.480 575.580 1391.600 ;
  LAYER metal1 ;
  RECT 572.040 1390.480 575.580 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 563.360 1390.480 566.900 1391.600 ;
  LAYER metal3 ;
  RECT 563.360 1390.480 566.900 1391.600 ;
  LAYER metal2 ;
  RECT 563.360 1390.480 566.900 1391.600 ;
  LAYER metal1 ;
  RECT 563.360 1390.480 566.900 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 554.680 1390.480 558.220 1391.600 ;
  LAYER metal3 ;
  RECT 554.680 1390.480 558.220 1391.600 ;
  LAYER metal2 ;
  RECT 554.680 1390.480 558.220 1391.600 ;
  LAYER metal1 ;
  RECT 554.680 1390.480 558.220 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 546.000 1390.480 549.540 1391.600 ;
  LAYER metal3 ;
  RECT 546.000 1390.480 549.540 1391.600 ;
  LAYER metal2 ;
  RECT 546.000 1390.480 549.540 1391.600 ;
  LAYER metal1 ;
  RECT 546.000 1390.480 549.540 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 537.320 1390.480 540.860 1391.600 ;
  LAYER metal3 ;
  RECT 537.320 1390.480 540.860 1391.600 ;
  LAYER metal2 ;
  RECT 537.320 1390.480 540.860 1391.600 ;
  LAYER metal1 ;
  RECT 537.320 1390.480 540.860 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 528.640 1390.480 532.180 1391.600 ;
  LAYER metal3 ;
  RECT 528.640 1390.480 532.180 1391.600 ;
  LAYER metal2 ;
  RECT 528.640 1390.480 532.180 1391.600 ;
  LAYER metal1 ;
  RECT 528.640 1390.480 532.180 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 485.240 1390.480 488.780 1391.600 ;
  LAYER metal3 ;
  RECT 485.240 1390.480 488.780 1391.600 ;
  LAYER metal2 ;
  RECT 485.240 1390.480 488.780 1391.600 ;
  LAYER metal1 ;
  RECT 485.240 1390.480 488.780 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 476.560 1390.480 480.100 1391.600 ;
  LAYER metal3 ;
  RECT 476.560 1390.480 480.100 1391.600 ;
  LAYER metal2 ;
  RECT 476.560 1390.480 480.100 1391.600 ;
  LAYER metal1 ;
  RECT 476.560 1390.480 480.100 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 467.880 1390.480 471.420 1391.600 ;
  LAYER metal3 ;
  RECT 467.880 1390.480 471.420 1391.600 ;
  LAYER metal2 ;
  RECT 467.880 1390.480 471.420 1391.600 ;
  LAYER metal1 ;
  RECT 467.880 1390.480 471.420 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 459.200 1390.480 462.740 1391.600 ;
  LAYER metal3 ;
  RECT 459.200 1390.480 462.740 1391.600 ;
  LAYER metal2 ;
  RECT 459.200 1390.480 462.740 1391.600 ;
  LAYER metal1 ;
  RECT 459.200 1390.480 462.740 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 450.520 1390.480 454.060 1391.600 ;
  LAYER metal3 ;
  RECT 450.520 1390.480 454.060 1391.600 ;
  LAYER metal2 ;
  RECT 450.520 1390.480 454.060 1391.600 ;
  LAYER metal1 ;
  RECT 450.520 1390.480 454.060 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 441.840 1390.480 445.380 1391.600 ;
  LAYER metal3 ;
  RECT 441.840 1390.480 445.380 1391.600 ;
  LAYER metal2 ;
  RECT 441.840 1390.480 445.380 1391.600 ;
  LAYER metal1 ;
  RECT 441.840 1390.480 445.380 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 398.440 1390.480 401.980 1391.600 ;
  LAYER metal3 ;
  RECT 398.440 1390.480 401.980 1391.600 ;
  LAYER metal2 ;
  RECT 398.440 1390.480 401.980 1391.600 ;
  LAYER metal1 ;
  RECT 398.440 1390.480 401.980 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 389.760 1390.480 393.300 1391.600 ;
  LAYER metal3 ;
  RECT 389.760 1390.480 393.300 1391.600 ;
  LAYER metal2 ;
  RECT 389.760 1390.480 393.300 1391.600 ;
  LAYER metal1 ;
  RECT 389.760 1390.480 393.300 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 381.080 1390.480 384.620 1391.600 ;
  LAYER metal3 ;
  RECT 381.080 1390.480 384.620 1391.600 ;
  LAYER metal2 ;
  RECT 381.080 1390.480 384.620 1391.600 ;
  LAYER metal1 ;
  RECT 381.080 1390.480 384.620 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 372.400 1390.480 375.940 1391.600 ;
  LAYER metal3 ;
  RECT 372.400 1390.480 375.940 1391.600 ;
  LAYER metal2 ;
  RECT 372.400 1390.480 375.940 1391.600 ;
  LAYER metal1 ;
  RECT 372.400 1390.480 375.940 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 363.720 1390.480 367.260 1391.600 ;
  LAYER metal3 ;
  RECT 363.720 1390.480 367.260 1391.600 ;
  LAYER metal2 ;
  RECT 363.720 1390.480 367.260 1391.600 ;
  LAYER metal1 ;
  RECT 363.720 1390.480 367.260 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 355.040 1390.480 358.580 1391.600 ;
  LAYER metal3 ;
  RECT 355.040 1390.480 358.580 1391.600 ;
  LAYER metal2 ;
  RECT 355.040 1390.480 358.580 1391.600 ;
  LAYER metal1 ;
  RECT 355.040 1390.480 358.580 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 311.640 1390.480 315.180 1391.600 ;
  LAYER metal3 ;
  RECT 311.640 1390.480 315.180 1391.600 ;
  LAYER metal2 ;
  RECT 311.640 1390.480 315.180 1391.600 ;
  LAYER metal1 ;
  RECT 311.640 1390.480 315.180 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 302.960 1390.480 306.500 1391.600 ;
  LAYER metal3 ;
  RECT 302.960 1390.480 306.500 1391.600 ;
  LAYER metal2 ;
  RECT 302.960 1390.480 306.500 1391.600 ;
  LAYER metal1 ;
  RECT 302.960 1390.480 306.500 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 294.280 1390.480 297.820 1391.600 ;
  LAYER metal3 ;
  RECT 294.280 1390.480 297.820 1391.600 ;
  LAYER metal2 ;
  RECT 294.280 1390.480 297.820 1391.600 ;
  LAYER metal1 ;
  RECT 294.280 1390.480 297.820 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 285.600 1390.480 289.140 1391.600 ;
  LAYER metal3 ;
  RECT 285.600 1390.480 289.140 1391.600 ;
  LAYER metal2 ;
  RECT 285.600 1390.480 289.140 1391.600 ;
  LAYER metal1 ;
  RECT 285.600 1390.480 289.140 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 276.920 1390.480 280.460 1391.600 ;
  LAYER metal3 ;
  RECT 276.920 1390.480 280.460 1391.600 ;
  LAYER metal2 ;
  RECT 276.920 1390.480 280.460 1391.600 ;
  LAYER metal1 ;
  RECT 276.920 1390.480 280.460 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 268.240 1390.480 271.780 1391.600 ;
  LAYER metal3 ;
  RECT 268.240 1390.480 271.780 1391.600 ;
  LAYER metal2 ;
  RECT 268.240 1390.480 271.780 1391.600 ;
  LAYER metal1 ;
  RECT 268.240 1390.480 271.780 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 224.840 1390.480 228.380 1391.600 ;
  LAYER metal3 ;
  RECT 224.840 1390.480 228.380 1391.600 ;
  LAYER metal2 ;
  RECT 224.840 1390.480 228.380 1391.600 ;
  LAYER metal1 ;
  RECT 224.840 1390.480 228.380 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 216.160 1390.480 219.700 1391.600 ;
  LAYER metal3 ;
  RECT 216.160 1390.480 219.700 1391.600 ;
  LAYER metal2 ;
  RECT 216.160 1390.480 219.700 1391.600 ;
  LAYER metal1 ;
  RECT 216.160 1390.480 219.700 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 207.480 1390.480 211.020 1391.600 ;
  LAYER metal3 ;
  RECT 207.480 1390.480 211.020 1391.600 ;
  LAYER metal2 ;
  RECT 207.480 1390.480 211.020 1391.600 ;
  LAYER metal1 ;
  RECT 207.480 1390.480 211.020 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.800 1390.480 202.340 1391.600 ;
  LAYER metal3 ;
  RECT 198.800 1390.480 202.340 1391.600 ;
  LAYER metal2 ;
  RECT 198.800 1390.480 202.340 1391.600 ;
  LAYER metal1 ;
  RECT 198.800 1390.480 202.340 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.120 1390.480 193.660 1391.600 ;
  LAYER metal3 ;
  RECT 190.120 1390.480 193.660 1391.600 ;
  LAYER metal2 ;
  RECT 190.120 1390.480 193.660 1391.600 ;
  LAYER metal1 ;
  RECT 190.120 1390.480 193.660 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 181.440 1390.480 184.980 1391.600 ;
  LAYER metal3 ;
  RECT 181.440 1390.480 184.980 1391.600 ;
  LAYER metal2 ;
  RECT 181.440 1390.480 184.980 1391.600 ;
  LAYER metal1 ;
  RECT 181.440 1390.480 184.980 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 138.040 1390.480 141.580 1391.600 ;
  LAYER metal3 ;
  RECT 138.040 1390.480 141.580 1391.600 ;
  LAYER metal2 ;
  RECT 138.040 1390.480 141.580 1391.600 ;
  LAYER metal1 ;
  RECT 138.040 1390.480 141.580 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 129.360 1390.480 132.900 1391.600 ;
  LAYER metal3 ;
  RECT 129.360 1390.480 132.900 1391.600 ;
  LAYER metal2 ;
  RECT 129.360 1390.480 132.900 1391.600 ;
  LAYER metal1 ;
  RECT 129.360 1390.480 132.900 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 120.680 1390.480 124.220 1391.600 ;
  LAYER metal3 ;
  RECT 120.680 1390.480 124.220 1391.600 ;
  LAYER metal2 ;
  RECT 120.680 1390.480 124.220 1391.600 ;
  LAYER metal1 ;
  RECT 120.680 1390.480 124.220 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 112.000 1390.480 115.540 1391.600 ;
  LAYER metal3 ;
  RECT 112.000 1390.480 115.540 1391.600 ;
  LAYER metal2 ;
  RECT 112.000 1390.480 115.540 1391.600 ;
  LAYER metal1 ;
  RECT 112.000 1390.480 115.540 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 103.320 1390.480 106.860 1391.600 ;
  LAYER metal3 ;
  RECT 103.320 1390.480 106.860 1391.600 ;
  LAYER metal2 ;
  RECT 103.320 1390.480 106.860 1391.600 ;
  LAYER metal1 ;
  RECT 103.320 1390.480 106.860 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 94.640 1390.480 98.180 1391.600 ;
  LAYER metal3 ;
  RECT 94.640 1390.480 98.180 1391.600 ;
  LAYER metal2 ;
  RECT 94.640 1390.480 98.180 1391.600 ;
  LAYER metal1 ;
  RECT 94.640 1390.480 98.180 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 51.240 1390.480 54.780 1391.600 ;
  LAYER metal3 ;
  RECT 51.240 1390.480 54.780 1391.600 ;
  LAYER metal2 ;
  RECT 51.240 1390.480 54.780 1391.600 ;
  LAYER metal1 ;
  RECT 51.240 1390.480 54.780 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 42.560 1390.480 46.100 1391.600 ;
  LAYER metal3 ;
  RECT 42.560 1390.480 46.100 1391.600 ;
  LAYER metal2 ;
  RECT 42.560 1390.480 46.100 1391.600 ;
  LAYER metal1 ;
  RECT 42.560 1390.480 46.100 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.880 1390.480 37.420 1391.600 ;
  LAYER metal3 ;
  RECT 33.880 1390.480 37.420 1391.600 ;
  LAYER metal2 ;
  RECT 33.880 1390.480 37.420 1391.600 ;
  LAYER metal1 ;
  RECT 33.880 1390.480 37.420 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.200 1390.480 28.740 1391.600 ;
  LAYER metal3 ;
  RECT 25.200 1390.480 28.740 1391.600 ;
  LAYER metal2 ;
  RECT 25.200 1390.480 28.740 1391.600 ;
  LAYER metal1 ;
  RECT 25.200 1390.480 28.740 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 16.520 1390.480 20.060 1391.600 ;
  LAYER metal3 ;
  RECT 16.520 1390.480 20.060 1391.600 ;
  LAYER metal2 ;
  RECT 16.520 1390.480 20.060 1391.600 ;
  LAYER metal1 ;
  RECT 16.520 1390.480 20.060 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.840 1390.480 11.380 1391.600 ;
  LAYER metal3 ;
  RECT 7.840 1390.480 11.380 1391.600 ;
  LAYER metal2 ;
  RECT 7.840 1390.480 11.380 1391.600 ;
  LAYER metal1 ;
  RECT 7.840 1390.480 11.380 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1908.760 0.000 1912.300 1.120 ;
  LAYER metal3 ;
  RECT 1908.760 0.000 1912.300 1.120 ;
  LAYER metal2 ;
  RECT 1908.760 0.000 1912.300 1.120 ;
  LAYER metal1 ;
  RECT 1908.760 0.000 1912.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1865.360 0.000 1868.900 1.120 ;
  LAYER metal3 ;
  RECT 1865.360 0.000 1868.900 1.120 ;
  LAYER metal2 ;
  RECT 1865.360 0.000 1868.900 1.120 ;
  LAYER metal1 ;
  RECT 1865.360 0.000 1868.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1856.680 0.000 1860.220 1.120 ;
  LAYER metal3 ;
  RECT 1856.680 0.000 1860.220 1.120 ;
  LAYER metal2 ;
  RECT 1856.680 0.000 1860.220 1.120 ;
  LAYER metal1 ;
  RECT 1856.680 0.000 1860.220 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1848.000 0.000 1851.540 1.120 ;
  LAYER metal3 ;
  RECT 1848.000 0.000 1851.540 1.120 ;
  LAYER metal2 ;
  RECT 1848.000 0.000 1851.540 1.120 ;
  LAYER metal1 ;
  RECT 1848.000 0.000 1851.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1839.320 0.000 1842.860 1.120 ;
  LAYER metal3 ;
  RECT 1839.320 0.000 1842.860 1.120 ;
  LAYER metal2 ;
  RECT 1839.320 0.000 1842.860 1.120 ;
  LAYER metal1 ;
  RECT 1839.320 0.000 1842.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1830.640 0.000 1834.180 1.120 ;
  LAYER metal3 ;
  RECT 1830.640 0.000 1834.180 1.120 ;
  LAYER metal2 ;
  RECT 1830.640 0.000 1834.180 1.120 ;
  LAYER metal1 ;
  RECT 1830.640 0.000 1834.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
  LAYER metal3 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
  LAYER metal2 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
  LAYER metal1 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1761.200 0.000 1764.740 1.120 ;
  LAYER metal3 ;
  RECT 1761.200 0.000 1764.740 1.120 ;
  LAYER metal2 ;
  RECT 1761.200 0.000 1764.740 1.120 ;
  LAYER metal1 ;
  RECT 1761.200 0.000 1764.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1752.520 0.000 1756.060 1.120 ;
  LAYER metal3 ;
  RECT 1752.520 0.000 1756.060 1.120 ;
  LAYER metal2 ;
  RECT 1752.520 0.000 1756.060 1.120 ;
  LAYER metal1 ;
  RECT 1752.520 0.000 1756.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1743.840 0.000 1747.380 1.120 ;
  LAYER metal3 ;
  RECT 1743.840 0.000 1747.380 1.120 ;
  LAYER metal2 ;
  RECT 1743.840 0.000 1747.380 1.120 ;
  LAYER metal1 ;
  RECT 1743.840 0.000 1747.380 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1735.160 0.000 1738.700 1.120 ;
  LAYER metal3 ;
  RECT 1735.160 0.000 1738.700 1.120 ;
  LAYER metal2 ;
  RECT 1735.160 0.000 1738.700 1.120 ;
  LAYER metal1 ;
  RECT 1735.160 0.000 1738.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1726.480 0.000 1730.020 1.120 ;
  LAYER metal3 ;
  RECT 1726.480 0.000 1730.020 1.120 ;
  LAYER metal2 ;
  RECT 1726.480 0.000 1730.020 1.120 ;
  LAYER metal1 ;
  RECT 1726.480 0.000 1730.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1717.800 0.000 1721.340 1.120 ;
  LAYER metal3 ;
  RECT 1717.800 0.000 1721.340 1.120 ;
  LAYER metal2 ;
  RECT 1717.800 0.000 1721.340 1.120 ;
  LAYER metal1 ;
  RECT 1717.800 0.000 1721.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1657.040 0.000 1660.580 1.120 ;
  LAYER metal3 ;
  RECT 1657.040 0.000 1660.580 1.120 ;
  LAYER metal2 ;
  RECT 1657.040 0.000 1660.580 1.120 ;
  LAYER metal1 ;
  RECT 1657.040 0.000 1660.580 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1648.360 0.000 1651.900 1.120 ;
  LAYER metal3 ;
  RECT 1648.360 0.000 1651.900 1.120 ;
  LAYER metal2 ;
  RECT 1648.360 0.000 1651.900 1.120 ;
  LAYER metal1 ;
  RECT 1648.360 0.000 1651.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1639.680 0.000 1643.220 1.120 ;
  LAYER metal3 ;
  RECT 1639.680 0.000 1643.220 1.120 ;
  LAYER metal2 ;
  RECT 1639.680 0.000 1643.220 1.120 ;
  LAYER metal1 ;
  RECT 1639.680 0.000 1643.220 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1631.000 0.000 1634.540 1.120 ;
  LAYER metal3 ;
  RECT 1631.000 0.000 1634.540 1.120 ;
  LAYER metal2 ;
  RECT 1631.000 0.000 1634.540 1.120 ;
  LAYER metal1 ;
  RECT 1631.000 0.000 1634.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1622.320 0.000 1625.860 1.120 ;
  LAYER metal3 ;
  RECT 1622.320 0.000 1625.860 1.120 ;
  LAYER metal2 ;
  RECT 1622.320 0.000 1625.860 1.120 ;
  LAYER metal1 ;
  RECT 1622.320 0.000 1625.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1613.640 0.000 1617.180 1.120 ;
  LAYER metal3 ;
  RECT 1613.640 0.000 1617.180 1.120 ;
  LAYER metal2 ;
  RECT 1613.640 0.000 1617.180 1.120 ;
  LAYER metal1 ;
  RECT 1613.640 0.000 1617.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1552.260 0.000 1555.800 1.120 ;
  LAYER metal3 ;
  RECT 1552.260 0.000 1555.800 1.120 ;
  LAYER metal2 ;
  RECT 1552.260 0.000 1555.800 1.120 ;
  LAYER metal1 ;
  RECT 1552.260 0.000 1555.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1543.580 0.000 1547.120 1.120 ;
  LAYER metal3 ;
  RECT 1543.580 0.000 1547.120 1.120 ;
  LAYER metal2 ;
  RECT 1543.580 0.000 1547.120 1.120 ;
  LAYER metal1 ;
  RECT 1543.580 0.000 1547.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1534.900 0.000 1538.440 1.120 ;
  LAYER metal3 ;
  RECT 1534.900 0.000 1538.440 1.120 ;
  LAYER metal2 ;
  RECT 1534.900 0.000 1538.440 1.120 ;
  LAYER metal1 ;
  RECT 1534.900 0.000 1538.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1526.220 0.000 1529.760 1.120 ;
  LAYER metal3 ;
  RECT 1526.220 0.000 1529.760 1.120 ;
  LAYER metal2 ;
  RECT 1526.220 0.000 1529.760 1.120 ;
  LAYER metal1 ;
  RECT 1526.220 0.000 1529.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1517.540 0.000 1521.080 1.120 ;
  LAYER metal3 ;
  RECT 1517.540 0.000 1521.080 1.120 ;
  LAYER metal2 ;
  RECT 1517.540 0.000 1521.080 1.120 ;
  LAYER metal1 ;
  RECT 1517.540 0.000 1521.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1508.860 0.000 1512.400 1.120 ;
  LAYER metal3 ;
  RECT 1508.860 0.000 1512.400 1.120 ;
  LAYER metal2 ;
  RECT 1508.860 0.000 1512.400 1.120 ;
  LAYER metal1 ;
  RECT 1508.860 0.000 1512.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1448.100 0.000 1451.640 1.120 ;
  LAYER metal3 ;
  RECT 1448.100 0.000 1451.640 1.120 ;
  LAYER metal2 ;
  RECT 1448.100 0.000 1451.640 1.120 ;
  LAYER metal1 ;
  RECT 1448.100 0.000 1451.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1439.420 0.000 1442.960 1.120 ;
  LAYER metal3 ;
  RECT 1439.420 0.000 1442.960 1.120 ;
  LAYER metal2 ;
  RECT 1439.420 0.000 1442.960 1.120 ;
  LAYER metal1 ;
  RECT 1439.420 0.000 1442.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1430.740 0.000 1434.280 1.120 ;
  LAYER metal3 ;
  RECT 1430.740 0.000 1434.280 1.120 ;
  LAYER metal2 ;
  RECT 1430.740 0.000 1434.280 1.120 ;
  LAYER metal1 ;
  RECT 1430.740 0.000 1434.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1422.060 0.000 1425.600 1.120 ;
  LAYER metal3 ;
  RECT 1422.060 0.000 1425.600 1.120 ;
  LAYER metal2 ;
  RECT 1422.060 0.000 1425.600 1.120 ;
  LAYER metal1 ;
  RECT 1422.060 0.000 1425.600 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1413.380 0.000 1416.920 1.120 ;
  LAYER metal3 ;
  RECT 1413.380 0.000 1416.920 1.120 ;
  LAYER metal2 ;
  RECT 1413.380 0.000 1416.920 1.120 ;
  LAYER metal1 ;
  RECT 1413.380 0.000 1416.920 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1404.700 0.000 1408.240 1.120 ;
  LAYER metal3 ;
  RECT 1404.700 0.000 1408.240 1.120 ;
  LAYER metal2 ;
  RECT 1404.700 0.000 1408.240 1.120 ;
  LAYER metal1 ;
  RECT 1404.700 0.000 1408.240 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1348.280 0.000 1351.820 1.120 ;
  LAYER metal3 ;
  RECT 1348.280 0.000 1351.820 1.120 ;
  LAYER metal2 ;
  RECT 1348.280 0.000 1351.820 1.120 ;
  LAYER metal1 ;
  RECT 1348.280 0.000 1351.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1335.260 0.000 1338.800 1.120 ;
  LAYER metal3 ;
  RECT 1335.260 0.000 1338.800 1.120 ;
  LAYER metal2 ;
  RECT 1335.260 0.000 1338.800 1.120 ;
  LAYER metal1 ;
  RECT 1335.260 0.000 1338.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1326.580 0.000 1330.120 1.120 ;
  LAYER metal3 ;
  RECT 1326.580 0.000 1330.120 1.120 ;
  LAYER metal2 ;
  RECT 1326.580 0.000 1330.120 1.120 ;
  LAYER metal1 ;
  RECT 1326.580 0.000 1330.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1317.900 0.000 1321.440 1.120 ;
  LAYER metal3 ;
  RECT 1317.900 0.000 1321.440 1.120 ;
  LAYER metal2 ;
  RECT 1317.900 0.000 1321.440 1.120 ;
  LAYER metal1 ;
  RECT 1317.900 0.000 1321.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1309.220 0.000 1312.760 1.120 ;
  LAYER metal3 ;
  RECT 1309.220 0.000 1312.760 1.120 ;
  LAYER metal2 ;
  RECT 1309.220 0.000 1312.760 1.120 ;
  LAYER metal1 ;
  RECT 1309.220 0.000 1312.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1300.540 0.000 1304.080 1.120 ;
  LAYER metal3 ;
  RECT 1300.540 0.000 1304.080 1.120 ;
  LAYER metal2 ;
  RECT 1300.540 0.000 1304.080 1.120 ;
  LAYER metal1 ;
  RECT 1300.540 0.000 1304.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1257.140 0.000 1260.680 1.120 ;
  LAYER metal3 ;
  RECT 1257.140 0.000 1260.680 1.120 ;
  LAYER metal2 ;
  RECT 1257.140 0.000 1260.680 1.120 ;
  LAYER metal1 ;
  RECT 1257.140 0.000 1260.680 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1235.440 0.000 1238.980 1.120 ;
  LAYER metal3 ;
  RECT 1235.440 0.000 1238.980 1.120 ;
  LAYER metal2 ;
  RECT 1235.440 0.000 1238.980 1.120 ;
  LAYER metal1 ;
  RECT 1235.440 0.000 1238.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1221.800 0.000 1225.340 1.120 ;
  LAYER metal3 ;
  RECT 1221.800 0.000 1225.340 1.120 ;
  LAYER metal2 ;
  RECT 1221.800 0.000 1225.340 1.120 ;
  LAYER metal1 ;
  RECT 1221.800 0.000 1225.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1213.120 0.000 1216.660 1.120 ;
  LAYER metal3 ;
  RECT 1213.120 0.000 1216.660 1.120 ;
  LAYER metal2 ;
  RECT 1213.120 0.000 1216.660 1.120 ;
  LAYER metal1 ;
  RECT 1213.120 0.000 1216.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1204.440 0.000 1207.980 1.120 ;
  LAYER metal3 ;
  RECT 1204.440 0.000 1207.980 1.120 ;
  LAYER metal2 ;
  RECT 1204.440 0.000 1207.980 1.120 ;
  LAYER metal1 ;
  RECT 1204.440 0.000 1207.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1195.760 0.000 1199.300 1.120 ;
  LAYER metal3 ;
  RECT 1195.760 0.000 1199.300 1.120 ;
  LAYER metal2 ;
  RECT 1195.760 0.000 1199.300 1.120 ;
  LAYER metal1 ;
  RECT 1195.760 0.000 1199.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1152.360 0.000 1155.900 1.120 ;
  LAYER metal3 ;
  RECT 1152.360 0.000 1155.900 1.120 ;
  LAYER metal2 ;
  RECT 1152.360 0.000 1155.900 1.120 ;
  LAYER metal1 ;
  RECT 1152.360 0.000 1155.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal3 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal2 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal1 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1121.980 0.000 1125.520 1.120 ;
  LAYER metal3 ;
  RECT 1121.980 0.000 1125.520 1.120 ;
  LAYER metal2 ;
  RECT 1121.980 0.000 1125.520 1.120 ;
  LAYER metal1 ;
  RECT 1121.980 0.000 1125.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1108.960 0.000 1112.500 1.120 ;
  LAYER metal3 ;
  RECT 1108.960 0.000 1112.500 1.120 ;
  LAYER metal2 ;
  RECT 1108.960 0.000 1112.500 1.120 ;
  LAYER metal1 ;
  RECT 1108.960 0.000 1112.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1100.280 0.000 1103.820 1.120 ;
  LAYER metal3 ;
  RECT 1100.280 0.000 1103.820 1.120 ;
  LAYER metal2 ;
  RECT 1100.280 0.000 1103.820 1.120 ;
  LAYER metal1 ;
  RECT 1100.280 0.000 1103.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1091.600 0.000 1095.140 1.120 ;
  LAYER metal3 ;
  RECT 1091.600 0.000 1095.140 1.120 ;
  LAYER metal2 ;
  RECT 1091.600 0.000 1095.140 1.120 ;
  LAYER metal1 ;
  RECT 1091.600 0.000 1095.140 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1048.200 0.000 1051.740 1.120 ;
  LAYER metal3 ;
  RECT 1048.200 0.000 1051.740 1.120 ;
  LAYER metal2 ;
  RECT 1048.200 0.000 1051.740 1.120 ;
  LAYER metal1 ;
  RECT 1048.200 0.000 1051.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1039.520 0.000 1043.060 1.120 ;
  LAYER metal3 ;
  RECT 1039.520 0.000 1043.060 1.120 ;
  LAYER metal2 ;
  RECT 1039.520 0.000 1043.060 1.120 ;
  LAYER metal1 ;
  RECT 1039.520 0.000 1043.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1030.840 0.000 1034.380 1.120 ;
  LAYER metal3 ;
  RECT 1030.840 0.000 1034.380 1.120 ;
  LAYER metal2 ;
  RECT 1030.840 0.000 1034.380 1.120 ;
  LAYER metal1 ;
  RECT 1030.840 0.000 1034.380 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1009.140 0.000 1012.680 1.120 ;
  LAYER metal3 ;
  RECT 1009.140 0.000 1012.680 1.120 ;
  LAYER metal2 ;
  RECT 1009.140 0.000 1012.680 1.120 ;
  LAYER metal1 ;
  RECT 1009.140 0.000 1012.680 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 977.520 0.000 981.060 1.120 ;
  LAYER metal3 ;
  RECT 977.520 0.000 981.060 1.120 ;
  LAYER metal2 ;
  RECT 977.520 0.000 981.060 1.120 ;
  LAYER metal1 ;
  RECT 977.520 0.000 981.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 956.440 0.000 959.980 1.120 ;
  LAYER metal3 ;
  RECT 956.440 0.000 959.980 1.120 ;
  LAYER metal2 ;
  RECT 956.440 0.000 959.980 1.120 ;
  LAYER metal1 ;
  RECT 956.440 0.000 959.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER metal3 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER metal2 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER metal1 ;
  RECT 887.620 0.000 891.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 878.940 0.000 882.480 1.120 ;
  LAYER metal3 ;
  RECT 878.940 0.000 882.480 1.120 ;
  LAYER metal2 ;
  RECT 878.940 0.000 882.480 1.120 ;
  LAYER metal1 ;
  RECT 878.940 0.000 882.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 870.260 0.000 873.800 1.120 ;
  LAYER metal3 ;
  RECT 870.260 0.000 873.800 1.120 ;
  LAYER metal2 ;
  RECT 870.260 0.000 873.800 1.120 ;
  LAYER metal1 ;
  RECT 870.260 0.000 873.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal3 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal2 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal1 ;
  RECT 861.580 0.000 865.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 852.900 0.000 856.440 1.120 ;
  LAYER metal3 ;
  RECT 852.900 0.000 856.440 1.120 ;
  LAYER metal2 ;
  RECT 852.900 0.000 856.440 1.120 ;
  LAYER metal1 ;
  RECT 852.900 0.000 856.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 844.220 0.000 847.760 1.120 ;
  LAYER metal3 ;
  RECT 844.220 0.000 847.760 1.120 ;
  LAYER metal2 ;
  RECT 844.220 0.000 847.760 1.120 ;
  LAYER metal1 ;
  RECT 844.220 0.000 847.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 783.460 0.000 787.000 1.120 ;
  LAYER metal3 ;
  RECT 783.460 0.000 787.000 1.120 ;
  LAYER metal2 ;
  RECT 783.460 0.000 787.000 1.120 ;
  LAYER metal1 ;
  RECT 783.460 0.000 787.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 774.780 0.000 778.320 1.120 ;
  LAYER metal3 ;
  RECT 774.780 0.000 778.320 1.120 ;
  LAYER metal2 ;
  RECT 774.780 0.000 778.320 1.120 ;
  LAYER metal1 ;
  RECT 774.780 0.000 778.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 766.100 0.000 769.640 1.120 ;
  LAYER metal3 ;
  RECT 766.100 0.000 769.640 1.120 ;
  LAYER metal2 ;
  RECT 766.100 0.000 769.640 1.120 ;
  LAYER metal1 ;
  RECT 766.100 0.000 769.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 757.420 0.000 760.960 1.120 ;
  LAYER metal3 ;
  RECT 757.420 0.000 760.960 1.120 ;
  LAYER metal2 ;
  RECT 757.420 0.000 760.960 1.120 ;
  LAYER metal1 ;
  RECT 757.420 0.000 760.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 748.740 0.000 752.280 1.120 ;
  LAYER metal3 ;
  RECT 748.740 0.000 752.280 1.120 ;
  LAYER metal2 ;
  RECT 748.740 0.000 752.280 1.120 ;
  LAYER metal1 ;
  RECT 748.740 0.000 752.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 740.060 0.000 743.600 1.120 ;
  LAYER metal3 ;
  RECT 740.060 0.000 743.600 1.120 ;
  LAYER metal2 ;
  RECT 740.060 0.000 743.600 1.120 ;
  LAYER metal1 ;
  RECT 740.060 0.000 743.600 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal3 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal2 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal1 ;
  RECT 678.680 0.000 682.220 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal3 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal2 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal1 ;
  RECT 670.000 0.000 673.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal3 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal2 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal1 ;
  RECT 661.320 0.000 664.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal3 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal2 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal1 ;
  RECT 652.640 0.000 656.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 643.960 0.000 647.500 1.120 ;
  LAYER metal3 ;
  RECT 643.960 0.000 647.500 1.120 ;
  LAYER metal2 ;
  RECT 643.960 0.000 647.500 1.120 ;
  LAYER metal1 ;
  RECT 643.960 0.000 647.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 635.280 0.000 638.820 1.120 ;
  LAYER metal3 ;
  RECT 635.280 0.000 638.820 1.120 ;
  LAYER metal2 ;
  RECT 635.280 0.000 638.820 1.120 ;
  LAYER metal1 ;
  RECT 635.280 0.000 638.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal3 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal2 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal1 ;
  RECT 578.860 0.000 582.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal3 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal2 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal1 ;
  RECT 565.840 0.000 569.380 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal3 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal2 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal1 ;
  RECT 557.160 0.000 560.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 548.480 0.000 552.020 1.120 ;
  LAYER metal3 ;
  RECT 548.480 0.000 552.020 1.120 ;
  LAYER metal2 ;
  RECT 548.480 0.000 552.020 1.120 ;
  LAYER metal1 ;
  RECT 548.480 0.000 552.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 539.800 0.000 543.340 1.120 ;
  LAYER metal3 ;
  RECT 539.800 0.000 543.340 1.120 ;
  LAYER metal2 ;
  RECT 539.800 0.000 543.340 1.120 ;
  LAYER metal1 ;
  RECT 539.800 0.000 543.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 531.120 0.000 534.660 1.120 ;
  LAYER metal3 ;
  RECT 531.120 0.000 534.660 1.120 ;
  LAYER metal2 ;
  RECT 531.120 0.000 534.660 1.120 ;
  LAYER metal1 ;
  RECT 531.120 0.000 534.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER metal3 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER metal2 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER metal1 ;
  RECT 487.720 0.000 491.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER metal3 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER metal2 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER metal1 ;
  RECT 466.020 0.000 469.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER metal3 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER metal2 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER metal1 ;
  RECT 453.000 0.000 456.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER metal3 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER metal2 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER metal1 ;
  RECT 444.320 0.000 447.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal3 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal2 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal1 ;
  RECT 435.640 0.000 439.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 426.960 0.000 430.500 1.120 ;
  LAYER metal3 ;
  RECT 426.960 0.000 430.500 1.120 ;
  LAYER metal2 ;
  RECT 426.960 0.000 430.500 1.120 ;
  LAYER metal1 ;
  RECT 426.960 0.000 430.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 383.560 0.000 387.100 1.120 ;
  LAYER metal3 ;
  RECT 383.560 0.000 387.100 1.120 ;
  LAYER metal2 ;
  RECT 383.560 0.000 387.100 1.120 ;
  LAYER metal1 ;
  RECT 383.560 0.000 387.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 374.880 0.000 378.420 1.120 ;
  LAYER metal3 ;
  RECT 374.880 0.000 378.420 1.120 ;
  LAYER metal2 ;
  RECT 374.880 0.000 378.420 1.120 ;
  LAYER metal1 ;
  RECT 374.880 0.000 378.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER metal3 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER metal2 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER metal1 ;
  RECT 353.180 0.000 356.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal3 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal2 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal1 ;
  RECT 339.540 0.000 343.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER metal3 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER metal2 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER metal1 ;
  RECT 330.860 0.000 334.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 322.180 0.000 325.720 1.120 ;
  LAYER metal3 ;
  RECT 322.180 0.000 325.720 1.120 ;
  LAYER metal2 ;
  RECT 322.180 0.000 325.720 1.120 ;
  LAYER metal1 ;
  RECT 322.180 0.000 325.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER metal3 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER metal2 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER metal1 ;
  RECT 278.780 0.000 282.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal3 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal2 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal1 ;
  RECT 270.100 0.000 273.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal3 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal2 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal1 ;
  RECT 261.420 0.000 264.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal3 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal2 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal1 ;
  RECT 239.720 0.000 243.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 226.700 0.000 230.240 1.120 ;
  LAYER metal3 ;
  RECT 226.700 0.000 230.240 1.120 ;
  LAYER metal2 ;
  RECT 226.700 0.000 230.240 1.120 ;
  LAYER metal1 ;
  RECT 226.700 0.000 230.240 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 218.020 0.000 221.560 1.120 ;
  LAYER metal3 ;
  RECT 218.020 0.000 221.560 1.120 ;
  LAYER metal2 ;
  RECT 218.020 0.000 221.560 1.120 ;
  LAYER metal1 ;
  RECT 218.020 0.000 221.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 174.620 0.000 178.160 1.120 ;
  LAYER metal3 ;
  RECT 174.620 0.000 178.160 1.120 ;
  LAYER metal2 ;
  RECT 174.620 0.000 178.160 1.120 ;
  LAYER metal1 ;
  RECT 174.620 0.000 178.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 165.940 0.000 169.480 1.120 ;
  LAYER metal3 ;
  RECT 165.940 0.000 169.480 1.120 ;
  LAYER metal2 ;
  RECT 165.940 0.000 169.480 1.120 ;
  LAYER metal1 ;
  RECT 165.940 0.000 169.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 157.260 0.000 160.800 1.120 ;
  LAYER metal3 ;
  RECT 157.260 0.000 160.800 1.120 ;
  LAYER metal2 ;
  RECT 157.260 0.000 160.800 1.120 ;
  LAYER metal1 ;
  RECT 157.260 0.000 160.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER metal3 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER metal2 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER metal1 ;
  RECT 148.580 0.000 152.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER metal3 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER metal2 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER metal1 ;
  RECT 61.780 0.000 65.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER metal3 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER metal2 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER metal1 ;
  RECT 53.100 0.000 56.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER metal3 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER metal2 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER metal1 ;
  RECT 44.420 0.000 47.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 1919.020 1376.260 1920.140 1379.500 ;
  LAYER metal3 ;
  RECT 1919.020 1376.260 1920.140 1379.500 ;
  LAYER metal2 ;
  RECT 1919.020 1376.260 1920.140 1379.500 ;
  LAYER metal1 ;
  RECT 1919.020 1376.260 1920.140 1379.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1368.420 1920.140 1371.660 ;
  LAYER metal3 ;
  RECT 1919.020 1368.420 1920.140 1371.660 ;
  LAYER metal2 ;
  RECT 1919.020 1368.420 1920.140 1371.660 ;
  LAYER metal1 ;
  RECT 1919.020 1368.420 1920.140 1371.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1360.580 1920.140 1363.820 ;
  LAYER metal3 ;
  RECT 1919.020 1360.580 1920.140 1363.820 ;
  LAYER metal2 ;
  RECT 1919.020 1360.580 1920.140 1363.820 ;
  LAYER metal1 ;
  RECT 1919.020 1360.580 1920.140 1363.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1352.740 1920.140 1355.980 ;
  LAYER metal3 ;
  RECT 1919.020 1352.740 1920.140 1355.980 ;
  LAYER metal2 ;
  RECT 1919.020 1352.740 1920.140 1355.980 ;
  LAYER metal1 ;
  RECT 1919.020 1352.740 1920.140 1355.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1344.900 1920.140 1348.140 ;
  LAYER metal3 ;
  RECT 1919.020 1344.900 1920.140 1348.140 ;
  LAYER metal2 ;
  RECT 1919.020 1344.900 1920.140 1348.140 ;
  LAYER metal1 ;
  RECT 1919.020 1344.900 1920.140 1348.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1305.700 1920.140 1308.940 ;
  LAYER metal3 ;
  RECT 1919.020 1305.700 1920.140 1308.940 ;
  LAYER metal2 ;
  RECT 1919.020 1305.700 1920.140 1308.940 ;
  LAYER metal1 ;
  RECT 1919.020 1305.700 1920.140 1308.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1297.860 1920.140 1301.100 ;
  LAYER metal3 ;
  RECT 1919.020 1297.860 1920.140 1301.100 ;
  LAYER metal2 ;
  RECT 1919.020 1297.860 1920.140 1301.100 ;
  LAYER metal1 ;
  RECT 1919.020 1297.860 1920.140 1301.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1290.020 1920.140 1293.260 ;
  LAYER metal3 ;
  RECT 1919.020 1290.020 1920.140 1293.260 ;
  LAYER metal2 ;
  RECT 1919.020 1290.020 1920.140 1293.260 ;
  LAYER metal1 ;
  RECT 1919.020 1290.020 1920.140 1293.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1282.180 1920.140 1285.420 ;
  LAYER metal3 ;
  RECT 1919.020 1282.180 1920.140 1285.420 ;
  LAYER metal2 ;
  RECT 1919.020 1282.180 1920.140 1285.420 ;
  LAYER metal1 ;
  RECT 1919.020 1282.180 1920.140 1285.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1274.340 1920.140 1277.580 ;
  LAYER metal3 ;
  RECT 1919.020 1274.340 1920.140 1277.580 ;
  LAYER metal2 ;
  RECT 1919.020 1274.340 1920.140 1277.580 ;
  LAYER metal1 ;
  RECT 1919.020 1274.340 1920.140 1277.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1266.500 1920.140 1269.740 ;
  LAYER metal3 ;
  RECT 1919.020 1266.500 1920.140 1269.740 ;
  LAYER metal2 ;
  RECT 1919.020 1266.500 1920.140 1269.740 ;
  LAYER metal1 ;
  RECT 1919.020 1266.500 1920.140 1269.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1227.300 1920.140 1230.540 ;
  LAYER metal3 ;
  RECT 1919.020 1227.300 1920.140 1230.540 ;
  LAYER metal2 ;
  RECT 1919.020 1227.300 1920.140 1230.540 ;
  LAYER metal1 ;
  RECT 1919.020 1227.300 1920.140 1230.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1219.460 1920.140 1222.700 ;
  LAYER metal3 ;
  RECT 1919.020 1219.460 1920.140 1222.700 ;
  LAYER metal2 ;
  RECT 1919.020 1219.460 1920.140 1222.700 ;
  LAYER metal1 ;
  RECT 1919.020 1219.460 1920.140 1222.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1211.620 1920.140 1214.860 ;
  LAYER metal3 ;
  RECT 1919.020 1211.620 1920.140 1214.860 ;
  LAYER metal2 ;
  RECT 1919.020 1211.620 1920.140 1214.860 ;
  LAYER metal1 ;
  RECT 1919.020 1211.620 1920.140 1214.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1203.780 1920.140 1207.020 ;
  LAYER metal3 ;
  RECT 1919.020 1203.780 1920.140 1207.020 ;
  LAYER metal2 ;
  RECT 1919.020 1203.780 1920.140 1207.020 ;
  LAYER metal1 ;
  RECT 1919.020 1203.780 1920.140 1207.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1195.940 1920.140 1199.180 ;
  LAYER metal3 ;
  RECT 1919.020 1195.940 1920.140 1199.180 ;
  LAYER metal2 ;
  RECT 1919.020 1195.940 1920.140 1199.180 ;
  LAYER metal1 ;
  RECT 1919.020 1195.940 1920.140 1199.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1188.100 1920.140 1191.340 ;
  LAYER metal3 ;
  RECT 1919.020 1188.100 1920.140 1191.340 ;
  LAYER metal2 ;
  RECT 1919.020 1188.100 1920.140 1191.340 ;
  LAYER metal1 ;
  RECT 1919.020 1188.100 1920.140 1191.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1148.900 1920.140 1152.140 ;
  LAYER metal3 ;
  RECT 1919.020 1148.900 1920.140 1152.140 ;
  LAYER metal2 ;
  RECT 1919.020 1148.900 1920.140 1152.140 ;
  LAYER metal1 ;
  RECT 1919.020 1148.900 1920.140 1152.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1141.060 1920.140 1144.300 ;
  LAYER metal3 ;
  RECT 1919.020 1141.060 1920.140 1144.300 ;
  LAYER metal2 ;
  RECT 1919.020 1141.060 1920.140 1144.300 ;
  LAYER metal1 ;
  RECT 1919.020 1141.060 1920.140 1144.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1133.220 1920.140 1136.460 ;
  LAYER metal3 ;
  RECT 1919.020 1133.220 1920.140 1136.460 ;
  LAYER metal2 ;
  RECT 1919.020 1133.220 1920.140 1136.460 ;
  LAYER metal1 ;
  RECT 1919.020 1133.220 1920.140 1136.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1125.380 1920.140 1128.620 ;
  LAYER metal3 ;
  RECT 1919.020 1125.380 1920.140 1128.620 ;
  LAYER metal2 ;
  RECT 1919.020 1125.380 1920.140 1128.620 ;
  LAYER metal1 ;
  RECT 1919.020 1125.380 1920.140 1128.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1117.540 1920.140 1120.780 ;
  LAYER metal3 ;
  RECT 1919.020 1117.540 1920.140 1120.780 ;
  LAYER metal2 ;
  RECT 1919.020 1117.540 1920.140 1120.780 ;
  LAYER metal1 ;
  RECT 1919.020 1117.540 1920.140 1120.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1109.700 1920.140 1112.940 ;
  LAYER metal3 ;
  RECT 1919.020 1109.700 1920.140 1112.940 ;
  LAYER metal2 ;
  RECT 1919.020 1109.700 1920.140 1112.940 ;
  LAYER metal1 ;
  RECT 1919.020 1109.700 1920.140 1112.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1070.500 1920.140 1073.740 ;
  LAYER metal3 ;
  RECT 1919.020 1070.500 1920.140 1073.740 ;
  LAYER metal2 ;
  RECT 1919.020 1070.500 1920.140 1073.740 ;
  LAYER metal1 ;
  RECT 1919.020 1070.500 1920.140 1073.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1062.660 1920.140 1065.900 ;
  LAYER metal3 ;
  RECT 1919.020 1062.660 1920.140 1065.900 ;
  LAYER metal2 ;
  RECT 1919.020 1062.660 1920.140 1065.900 ;
  LAYER metal1 ;
  RECT 1919.020 1062.660 1920.140 1065.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1054.820 1920.140 1058.060 ;
  LAYER metal3 ;
  RECT 1919.020 1054.820 1920.140 1058.060 ;
  LAYER metal2 ;
  RECT 1919.020 1054.820 1920.140 1058.060 ;
  LAYER metal1 ;
  RECT 1919.020 1054.820 1920.140 1058.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1046.980 1920.140 1050.220 ;
  LAYER metal3 ;
  RECT 1919.020 1046.980 1920.140 1050.220 ;
  LAYER metal2 ;
  RECT 1919.020 1046.980 1920.140 1050.220 ;
  LAYER metal1 ;
  RECT 1919.020 1046.980 1920.140 1050.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1039.140 1920.140 1042.380 ;
  LAYER metal3 ;
  RECT 1919.020 1039.140 1920.140 1042.380 ;
  LAYER metal2 ;
  RECT 1919.020 1039.140 1920.140 1042.380 ;
  LAYER metal1 ;
  RECT 1919.020 1039.140 1920.140 1042.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 1031.300 1920.140 1034.540 ;
  LAYER metal3 ;
  RECT 1919.020 1031.300 1920.140 1034.540 ;
  LAYER metal2 ;
  RECT 1919.020 1031.300 1920.140 1034.540 ;
  LAYER metal1 ;
  RECT 1919.020 1031.300 1920.140 1034.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 992.100 1920.140 995.340 ;
  LAYER metal3 ;
  RECT 1919.020 992.100 1920.140 995.340 ;
  LAYER metal2 ;
  RECT 1919.020 992.100 1920.140 995.340 ;
  LAYER metal1 ;
  RECT 1919.020 992.100 1920.140 995.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 984.260 1920.140 987.500 ;
  LAYER metal3 ;
  RECT 1919.020 984.260 1920.140 987.500 ;
  LAYER metal2 ;
  RECT 1919.020 984.260 1920.140 987.500 ;
  LAYER metal1 ;
  RECT 1919.020 984.260 1920.140 987.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 976.420 1920.140 979.660 ;
  LAYER metal3 ;
  RECT 1919.020 976.420 1920.140 979.660 ;
  LAYER metal2 ;
  RECT 1919.020 976.420 1920.140 979.660 ;
  LAYER metal1 ;
  RECT 1919.020 976.420 1920.140 979.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 968.580 1920.140 971.820 ;
  LAYER metal3 ;
  RECT 1919.020 968.580 1920.140 971.820 ;
  LAYER metal2 ;
  RECT 1919.020 968.580 1920.140 971.820 ;
  LAYER metal1 ;
  RECT 1919.020 968.580 1920.140 971.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 960.740 1920.140 963.980 ;
  LAYER metal3 ;
  RECT 1919.020 960.740 1920.140 963.980 ;
  LAYER metal2 ;
  RECT 1919.020 960.740 1920.140 963.980 ;
  LAYER metal1 ;
  RECT 1919.020 960.740 1920.140 963.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 952.900 1920.140 956.140 ;
  LAYER metal3 ;
  RECT 1919.020 952.900 1920.140 956.140 ;
  LAYER metal2 ;
  RECT 1919.020 952.900 1920.140 956.140 ;
  LAYER metal1 ;
  RECT 1919.020 952.900 1920.140 956.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 913.700 1920.140 916.940 ;
  LAYER metal3 ;
  RECT 1919.020 913.700 1920.140 916.940 ;
  LAYER metal2 ;
  RECT 1919.020 913.700 1920.140 916.940 ;
  LAYER metal1 ;
  RECT 1919.020 913.700 1920.140 916.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 905.860 1920.140 909.100 ;
  LAYER metal3 ;
  RECT 1919.020 905.860 1920.140 909.100 ;
  LAYER metal2 ;
  RECT 1919.020 905.860 1920.140 909.100 ;
  LAYER metal1 ;
  RECT 1919.020 905.860 1920.140 909.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 898.020 1920.140 901.260 ;
  LAYER metal3 ;
  RECT 1919.020 898.020 1920.140 901.260 ;
  LAYER metal2 ;
  RECT 1919.020 898.020 1920.140 901.260 ;
  LAYER metal1 ;
  RECT 1919.020 898.020 1920.140 901.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 890.180 1920.140 893.420 ;
  LAYER metal3 ;
  RECT 1919.020 890.180 1920.140 893.420 ;
  LAYER metal2 ;
  RECT 1919.020 890.180 1920.140 893.420 ;
  LAYER metal1 ;
  RECT 1919.020 890.180 1920.140 893.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 882.340 1920.140 885.580 ;
  LAYER metal3 ;
  RECT 1919.020 882.340 1920.140 885.580 ;
  LAYER metal2 ;
  RECT 1919.020 882.340 1920.140 885.580 ;
  LAYER metal1 ;
  RECT 1919.020 882.340 1920.140 885.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 874.500 1920.140 877.740 ;
  LAYER metal3 ;
  RECT 1919.020 874.500 1920.140 877.740 ;
  LAYER metal2 ;
  RECT 1919.020 874.500 1920.140 877.740 ;
  LAYER metal1 ;
  RECT 1919.020 874.500 1920.140 877.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 835.300 1920.140 838.540 ;
  LAYER metal3 ;
  RECT 1919.020 835.300 1920.140 838.540 ;
  LAYER metal2 ;
  RECT 1919.020 835.300 1920.140 838.540 ;
  LAYER metal1 ;
  RECT 1919.020 835.300 1920.140 838.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 827.460 1920.140 830.700 ;
  LAYER metal3 ;
  RECT 1919.020 827.460 1920.140 830.700 ;
  LAYER metal2 ;
  RECT 1919.020 827.460 1920.140 830.700 ;
  LAYER metal1 ;
  RECT 1919.020 827.460 1920.140 830.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 819.620 1920.140 822.860 ;
  LAYER metal3 ;
  RECT 1919.020 819.620 1920.140 822.860 ;
  LAYER metal2 ;
  RECT 1919.020 819.620 1920.140 822.860 ;
  LAYER metal1 ;
  RECT 1919.020 819.620 1920.140 822.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 811.780 1920.140 815.020 ;
  LAYER metal3 ;
  RECT 1919.020 811.780 1920.140 815.020 ;
  LAYER metal2 ;
  RECT 1919.020 811.780 1920.140 815.020 ;
  LAYER metal1 ;
  RECT 1919.020 811.780 1920.140 815.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 803.940 1920.140 807.180 ;
  LAYER metal3 ;
  RECT 1919.020 803.940 1920.140 807.180 ;
  LAYER metal2 ;
  RECT 1919.020 803.940 1920.140 807.180 ;
  LAYER metal1 ;
  RECT 1919.020 803.940 1920.140 807.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 796.100 1920.140 799.340 ;
  LAYER metal3 ;
  RECT 1919.020 796.100 1920.140 799.340 ;
  LAYER metal2 ;
  RECT 1919.020 796.100 1920.140 799.340 ;
  LAYER metal1 ;
  RECT 1919.020 796.100 1920.140 799.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 756.900 1920.140 760.140 ;
  LAYER metal3 ;
  RECT 1919.020 756.900 1920.140 760.140 ;
  LAYER metal2 ;
  RECT 1919.020 756.900 1920.140 760.140 ;
  LAYER metal1 ;
  RECT 1919.020 756.900 1920.140 760.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 749.060 1920.140 752.300 ;
  LAYER metal3 ;
  RECT 1919.020 749.060 1920.140 752.300 ;
  LAYER metal2 ;
  RECT 1919.020 749.060 1920.140 752.300 ;
  LAYER metal1 ;
  RECT 1919.020 749.060 1920.140 752.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 741.220 1920.140 744.460 ;
  LAYER metal3 ;
  RECT 1919.020 741.220 1920.140 744.460 ;
  LAYER metal2 ;
  RECT 1919.020 741.220 1920.140 744.460 ;
  LAYER metal1 ;
  RECT 1919.020 741.220 1920.140 744.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 733.380 1920.140 736.620 ;
  LAYER metal3 ;
  RECT 1919.020 733.380 1920.140 736.620 ;
  LAYER metal2 ;
  RECT 1919.020 733.380 1920.140 736.620 ;
  LAYER metal1 ;
  RECT 1919.020 733.380 1920.140 736.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 725.540 1920.140 728.780 ;
  LAYER metal3 ;
  RECT 1919.020 725.540 1920.140 728.780 ;
  LAYER metal2 ;
  RECT 1919.020 725.540 1920.140 728.780 ;
  LAYER metal1 ;
  RECT 1919.020 725.540 1920.140 728.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 717.700 1920.140 720.940 ;
  LAYER metal3 ;
  RECT 1919.020 717.700 1920.140 720.940 ;
  LAYER metal2 ;
  RECT 1919.020 717.700 1920.140 720.940 ;
  LAYER metal1 ;
  RECT 1919.020 717.700 1920.140 720.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 678.500 1920.140 681.740 ;
  LAYER metal3 ;
  RECT 1919.020 678.500 1920.140 681.740 ;
  LAYER metal2 ;
  RECT 1919.020 678.500 1920.140 681.740 ;
  LAYER metal1 ;
  RECT 1919.020 678.500 1920.140 681.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 670.660 1920.140 673.900 ;
  LAYER metal3 ;
  RECT 1919.020 670.660 1920.140 673.900 ;
  LAYER metal2 ;
  RECT 1919.020 670.660 1920.140 673.900 ;
  LAYER metal1 ;
  RECT 1919.020 670.660 1920.140 673.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 662.820 1920.140 666.060 ;
  LAYER metal3 ;
  RECT 1919.020 662.820 1920.140 666.060 ;
  LAYER metal2 ;
  RECT 1919.020 662.820 1920.140 666.060 ;
  LAYER metal1 ;
  RECT 1919.020 662.820 1920.140 666.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 654.980 1920.140 658.220 ;
  LAYER metal3 ;
  RECT 1919.020 654.980 1920.140 658.220 ;
  LAYER metal2 ;
  RECT 1919.020 654.980 1920.140 658.220 ;
  LAYER metal1 ;
  RECT 1919.020 654.980 1920.140 658.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 647.140 1920.140 650.380 ;
  LAYER metal3 ;
  RECT 1919.020 647.140 1920.140 650.380 ;
  LAYER metal2 ;
  RECT 1919.020 647.140 1920.140 650.380 ;
  LAYER metal1 ;
  RECT 1919.020 647.140 1920.140 650.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 639.300 1920.140 642.540 ;
  LAYER metal3 ;
  RECT 1919.020 639.300 1920.140 642.540 ;
  LAYER metal2 ;
  RECT 1919.020 639.300 1920.140 642.540 ;
  LAYER metal1 ;
  RECT 1919.020 639.300 1920.140 642.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 600.100 1920.140 603.340 ;
  LAYER metal3 ;
  RECT 1919.020 600.100 1920.140 603.340 ;
  LAYER metal2 ;
  RECT 1919.020 600.100 1920.140 603.340 ;
  LAYER metal1 ;
  RECT 1919.020 600.100 1920.140 603.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 592.260 1920.140 595.500 ;
  LAYER metal3 ;
  RECT 1919.020 592.260 1920.140 595.500 ;
  LAYER metal2 ;
  RECT 1919.020 592.260 1920.140 595.500 ;
  LAYER metal1 ;
  RECT 1919.020 592.260 1920.140 595.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 584.420 1920.140 587.660 ;
  LAYER metal3 ;
  RECT 1919.020 584.420 1920.140 587.660 ;
  LAYER metal2 ;
  RECT 1919.020 584.420 1920.140 587.660 ;
  LAYER metal1 ;
  RECT 1919.020 584.420 1920.140 587.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 576.580 1920.140 579.820 ;
  LAYER metal3 ;
  RECT 1919.020 576.580 1920.140 579.820 ;
  LAYER metal2 ;
  RECT 1919.020 576.580 1920.140 579.820 ;
  LAYER metal1 ;
  RECT 1919.020 576.580 1920.140 579.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 568.740 1920.140 571.980 ;
  LAYER metal3 ;
  RECT 1919.020 568.740 1920.140 571.980 ;
  LAYER metal2 ;
  RECT 1919.020 568.740 1920.140 571.980 ;
  LAYER metal1 ;
  RECT 1919.020 568.740 1920.140 571.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 560.900 1920.140 564.140 ;
  LAYER metal3 ;
  RECT 1919.020 560.900 1920.140 564.140 ;
  LAYER metal2 ;
  RECT 1919.020 560.900 1920.140 564.140 ;
  LAYER metal1 ;
  RECT 1919.020 560.900 1920.140 564.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 521.700 1920.140 524.940 ;
  LAYER metal3 ;
  RECT 1919.020 521.700 1920.140 524.940 ;
  LAYER metal2 ;
  RECT 1919.020 521.700 1920.140 524.940 ;
  LAYER metal1 ;
  RECT 1919.020 521.700 1920.140 524.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 513.860 1920.140 517.100 ;
  LAYER metal3 ;
  RECT 1919.020 513.860 1920.140 517.100 ;
  LAYER metal2 ;
  RECT 1919.020 513.860 1920.140 517.100 ;
  LAYER metal1 ;
  RECT 1919.020 513.860 1920.140 517.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 506.020 1920.140 509.260 ;
  LAYER metal3 ;
  RECT 1919.020 506.020 1920.140 509.260 ;
  LAYER metal2 ;
  RECT 1919.020 506.020 1920.140 509.260 ;
  LAYER metal1 ;
  RECT 1919.020 506.020 1920.140 509.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 498.180 1920.140 501.420 ;
  LAYER metal3 ;
  RECT 1919.020 498.180 1920.140 501.420 ;
  LAYER metal2 ;
  RECT 1919.020 498.180 1920.140 501.420 ;
  LAYER metal1 ;
  RECT 1919.020 498.180 1920.140 501.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 490.340 1920.140 493.580 ;
  LAYER metal3 ;
  RECT 1919.020 490.340 1920.140 493.580 ;
  LAYER metal2 ;
  RECT 1919.020 490.340 1920.140 493.580 ;
  LAYER metal1 ;
  RECT 1919.020 490.340 1920.140 493.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 482.500 1920.140 485.740 ;
  LAYER metal3 ;
  RECT 1919.020 482.500 1920.140 485.740 ;
  LAYER metal2 ;
  RECT 1919.020 482.500 1920.140 485.740 ;
  LAYER metal1 ;
  RECT 1919.020 482.500 1920.140 485.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 443.300 1920.140 446.540 ;
  LAYER metal3 ;
  RECT 1919.020 443.300 1920.140 446.540 ;
  LAYER metal2 ;
  RECT 1919.020 443.300 1920.140 446.540 ;
  LAYER metal1 ;
  RECT 1919.020 443.300 1920.140 446.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 435.460 1920.140 438.700 ;
  LAYER metal3 ;
  RECT 1919.020 435.460 1920.140 438.700 ;
  LAYER metal2 ;
  RECT 1919.020 435.460 1920.140 438.700 ;
  LAYER metal1 ;
  RECT 1919.020 435.460 1920.140 438.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 427.620 1920.140 430.860 ;
  LAYER metal3 ;
  RECT 1919.020 427.620 1920.140 430.860 ;
  LAYER metal2 ;
  RECT 1919.020 427.620 1920.140 430.860 ;
  LAYER metal1 ;
  RECT 1919.020 427.620 1920.140 430.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 419.780 1920.140 423.020 ;
  LAYER metal3 ;
  RECT 1919.020 419.780 1920.140 423.020 ;
  LAYER metal2 ;
  RECT 1919.020 419.780 1920.140 423.020 ;
  LAYER metal1 ;
  RECT 1919.020 419.780 1920.140 423.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 411.940 1920.140 415.180 ;
  LAYER metal3 ;
  RECT 1919.020 411.940 1920.140 415.180 ;
  LAYER metal2 ;
  RECT 1919.020 411.940 1920.140 415.180 ;
  LAYER metal1 ;
  RECT 1919.020 411.940 1920.140 415.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 404.100 1920.140 407.340 ;
  LAYER metal3 ;
  RECT 1919.020 404.100 1920.140 407.340 ;
  LAYER metal2 ;
  RECT 1919.020 404.100 1920.140 407.340 ;
  LAYER metal1 ;
  RECT 1919.020 404.100 1920.140 407.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 364.900 1920.140 368.140 ;
  LAYER metal3 ;
  RECT 1919.020 364.900 1920.140 368.140 ;
  LAYER metal2 ;
  RECT 1919.020 364.900 1920.140 368.140 ;
  LAYER metal1 ;
  RECT 1919.020 364.900 1920.140 368.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 357.060 1920.140 360.300 ;
  LAYER metal3 ;
  RECT 1919.020 357.060 1920.140 360.300 ;
  LAYER metal2 ;
  RECT 1919.020 357.060 1920.140 360.300 ;
  LAYER metal1 ;
  RECT 1919.020 357.060 1920.140 360.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 349.220 1920.140 352.460 ;
  LAYER metal3 ;
  RECT 1919.020 349.220 1920.140 352.460 ;
  LAYER metal2 ;
  RECT 1919.020 349.220 1920.140 352.460 ;
  LAYER metal1 ;
  RECT 1919.020 349.220 1920.140 352.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 341.380 1920.140 344.620 ;
  LAYER metal3 ;
  RECT 1919.020 341.380 1920.140 344.620 ;
  LAYER metal2 ;
  RECT 1919.020 341.380 1920.140 344.620 ;
  LAYER metal1 ;
  RECT 1919.020 341.380 1920.140 344.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 333.540 1920.140 336.780 ;
  LAYER metal3 ;
  RECT 1919.020 333.540 1920.140 336.780 ;
  LAYER metal2 ;
  RECT 1919.020 333.540 1920.140 336.780 ;
  LAYER metal1 ;
  RECT 1919.020 333.540 1920.140 336.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 325.700 1920.140 328.940 ;
  LAYER metal3 ;
  RECT 1919.020 325.700 1920.140 328.940 ;
  LAYER metal2 ;
  RECT 1919.020 325.700 1920.140 328.940 ;
  LAYER metal1 ;
  RECT 1919.020 325.700 1920.140 328.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 286.500 1920.140 289.740 ;
  LAYER metal3 ;
  RECT 1919.020 286.500 1920.140 289.740 ;
  LAYER metal2 ;
  RECT 1919.020 286.500 1920.140 289.740 ;
  LAYER metal1 ;
  RECT 1919.020 286.500 1920.140 289.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 278.660 1920.140 281.900 ;
  LAYER metal3 ;
  RECT 1919.020 278.660 1920.140 281.900 ;
  LAYER metal2 ;
  RECT 1919.020 278.660 1920.140 281.900 ;
  LAYER metal1 ;
  RECT 1919.020 278.660 1920.140 281.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 270.820 1920.140 274.060 ;
  LAYER metal3 ;
  RECT 1919.020 270.820 1920.140 274.060 ;
  LAYER metal2 ;
  RECT 1919.020 270.820 1920.140 274.060 ;
  LAYER metal1 ;
  RECT 1919.020 270.820 1920.140 274.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 262.980 1920.140 266.220 ;
  LAYER metal3 ;
  RECT 1919.020 262.980 1920.140 266.220 ;
  LAYER metal2 ;
  RECT 1919.020 262.980 1920.140 266.220 ;
  LAYER metal1 ;
  RECT 1919.020 262.980 1920.140 266.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 255.140 1920.140 258.380 ;
  LAYER metal3 ;
  RECT 1919.020 255.140 1920.140 258.380 ;
  LAYER metal2 ;
  RECT 1919.020 255.140 1920.140 258.380 ;
  LAYER metal1 ;
  RECT 1919.020 255.140 1920.140 258.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 247.300 1920.140 250.540 ;
  LAYER metal3 ;
  RECT 1919.020 247.300 1920.140 250.540 ;
  LAYER metal2 ;
  RECT 1919.020 247.300 1920.140 250.540 ;
  LAYER metal1 ;
  RECT 1919.020 247.300 1920.140 250.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 208.100 1920.140 211.340 ;
  LAYER metal3 ;
  RECT 1919.020 208.100 1920.140 211.340 ;
  LAYER metal2 ;
  RECT 1919.020 208.100 1920.140 211.340 ;
  LAYER metal1 ;
  RECT 1919.020 208.100 1920.140 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 200.260 1920.140 203.500 ;
  LAYER metal3 ;
  RECT 1919.020 200.260 1920.140 203.500 ;
  LAYER metal2 ;
  RECT 1919.020 200.260 1920.140 203.500 ;
  LAYER metal1 ;
  RECT 1919.020 200.260 1920.140 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 192.420 1920.140 195.660 ;
  LAYER metal3 ;
  RECT 1919.020 192.420 1920.140 195.660 ;
  LAYER metal2 ;
  RECT 1919.020 192.420 1920.140 195.660 ;
  LAYER metal1 ;
  RECT 1919.020 192.420 1920.140 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 184.580 1920.140 187.820 ;
  LAYER metal3 ;
  RECT 1919.020 184.580 1920.140 187.820 ;
  LAYER metal2 ;
  RECT 1919.020 184.580 1920.140 187.820 ;
  LAYER metal1 ;
  RECT 1919.020 184.580 1920.140 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 176.740 1920.140 179.980 ;
  LAYER metal3 ;
  RECT 1919.020 176.740 1920.140 179.980 ;
  LAYER metal2 ;
  RECT 1919.020 176.740 1920.140 179.980 ;
  LAYER metal1 ;
  RECT 1919.020 176.740 1920.140 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 168.900 1920.140 172.140 ;
  LAYER metal3 ;
  RECT 1919.020 168.900 1920.140 172.140 ;
  LAYER metal2 ;
  RECT 1919.020 168.900 1920.140 172.140 ;
  LAYER metal1 ;
  RECT 1919.020 168.900 1920.140 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 129.700 1920.140 132.940 ;
  LAYER metal3 ;
  RECT 1919.020 129.700 1920.140 132.940 ;
  LAYER metal2 ;
  RECT 1919.020 129.700 1920.140 132.940 ;
  LAYER metal1 ;
  RECT 1919.020 129.700 1920.140 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 121.860 1920.140 125.100 ;
  LAYER metal3 ;
  RECT 1919.020 121.860 1920.140 125.100 ;
  LAYER metal2 ;
  RECT 1919.020 121.860 1920.140 125.100 ;
  LAYER metal1 ;
  RECT 1919.020 121.860 1920.140 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 114.020 1920.140 117.260 ;
  LAYER metal3 ;
  RECT 1919.020 114.020 1920.140 117.260 ;
  LAYER metal2 ;
  RECT 1919.020 114.020 1920.140 117.260 ;
  LAYER metal1 ;
  RECT 1919.020 114.020 1920.140 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 106.180 1920.140 109.420 ;
  LAYER metal3 ;
  RECT 1919.020 106.180 1920.140 109.420 ;
  LAYER metal2 ;
  RECT 1919.020 106.180 1920.140 109.420 ;
  LAYER metal1 ;
  RECT 1919.020 106.180 1920.140 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 98.340 1920.140 101.580 ;
  LAYER metal3 ;
  RECT 1919.020 98.340 1920.140 101.580 ;
  LAYER metal2 ;
  RECT 1919.020 98.340 1920.140 101.580 ;
  LAYER metal1 ;
  RECT 1919.020 98.340 1920.140 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 90.500 1920.140 93.740 ;
  LAYER metal3 ;
  RECT 1919.020 90.500 1920.140 93.740 ;
  LAYER metal2 ;
  RECT 1919.020 90.500 1920.140 93.740 ;
  LAYER metal1 ;
  RECT 1919.020 90.500 1920.140 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 51.300 1920.140 54.540 ;
  LAYER metal3 ;
  RECT 1919.020 51.300 1920.140 54.540 ;
  LAYER metal2 ;
  RECT 1919.020 51.300 1920.140 54.540 ;
  LAYER metal1 ;
  RECT 1919.020 51.300 1920.140 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 43.460 1920.140 46.700 ;
  LAYER metal3 ;
  RECT 1919.020 43.460 1920.140 46.700 ;
  LAYER metal2 ;
  RECT 1919.020 43.460 1920.140 46.700 ;
  LAYER metal1 ;
  RECT 1919.020 43.460 1920.140 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 35.620 1920.140 38.860 ;
  LAYER metal3 ;
  RECT 1919.020 35.620 1920.140 38.860 ;
  LAYER metal2 ;
  RECT 1919.020 35.620 1920.140 38.860 ;
  LAYER metal1 ;
  RECT 1919.020 35.620 1920.140 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 27.780 1920.140 31.020 ;
  LAYER metal3 ;
  RECT 1919.020 27.780 1920.140 31.020 ;
  LAYER metal2 ;
  RECT 1919.020 27.780 1920.140 31.020 ;
  LAYER metal1 ;
  RECT 1919.020 27.780 1920.140 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 19.940 1920.140 23.180 ;
  LAYER metal3 ;
  RECT 1919.020 19.940 1920.140 23.180 ;
  LAYER metal2 ;
  RECT 1919.020 19.940 1920.140 23.180 ;
  LAYER metal1 ;
  RECT 1919.020 19.940 1920.140 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1919.020 12.100 1920.140 15.340 ;
  LAYER metal3 ;
  RECT 1919.020 12.100 1920.140 15.340 ;
  LAYER metal2 ;
  RECT 1919.020 12.100 1920.140 15.340 ;
  LAYER metal1 ;
  RECT 1919.020 12.100 1920.140 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1376.260 1.120 1379.500 ;
  LAYER metal3 ;
  RECT 0.000 1376.260 1.120 1379.500 ;
  LAYER metal2 ;
  RECT 0.000 1376.260 1.120 1379.500 ;
  LAYER metal1 ;
  RECT 0.000 1376.260 1.120 1379.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1368.420 1.120 1371.660 ;
  LAYER metal3 ;
  RECT 0.000 1368.420 1.120 1371.660 ;
  LAYER metal2 ;
  RECT 0.000 1368.420 1.120 1371.660 ;
  LAYER metal1 ;
  RECT 0.000 1368.420 1.120 1371.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1360.580 1.120 1363.820 ;
  LAYER metal3 ;
  RECT 0.000 1360.580 1.120 1363.820 ;
  LAYER metal2 ;
  RECT 0.000 1360.580 1.120 1363.820 ;
  LAYER metal1 ;
  RECT 0.000 1360.580 1.120 1363.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1352.740 1.120 1355.980 ;
  LAYER metal3 ;
  RECT 0.000 1352.740 1.120 1355.980 ;
  LAYER metal2 ;
  RECT 0.000 1352.740 1.120 1355.980 ;
  LAYER metal1 ;
  RECT 0.000 1352.740 1.120 1355.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1344.900 1.120 1348.140 ;
  LAYER metal3 ;
  RECT 0.000 1344.900 1.120 1348.140 ;
  LAYER metal2 ;
  RECT 0.000 1344.900 1.120 1348.140 ;
  LAYER metal1 ;
  RECT 0.000 1344.900 1.120 1348.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1305.700 1.120 1308.940 ;
  LAYER metal3 ;
  RECT 0.000 1305.700 1.120 1308.940 ;
  LAYER metal2 ;
  RECT 0.000 1305.700 1.120 1308.940 ;
  LAYER metal1 ;
  RECT 0.000 1305.700 1.120 1308.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1297.860 1.120 1301.100 ;
  LAYER metal3 ;
  RECT 0.000 1297.860 1.120 1301.100 ;
  LAYER metal2 ;
  RECT 0.000 1297.860 1.120 1301.100 ;
  LAYER metal1 ;
  RECT 0.000 1297.860 1.120 1301.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1290.020 1.120 1293.260 ;
  LAYER metal3 ;
  RECT 0.000 1290.020 1.120 1293.260 ;
  LAYER metal2 ;
  RECT 0.000 1290.020 1.120 1293.260 ;
  LAYER metal1 ;
  RECT 0.000 1290.020 1.120 1293.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1282.180 1.120 1285.420 ;
  LAYER metal3 ;
  RECT 0.000 1282.180 1.120 1285.420 ;
  LAYER metal2 ;
  RECT 0.000 1282.180 1.120 1285.420 ;
  LAYER metal1 ;
  RECT 0.000 1282.180 1.120 1285.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1274.340 1.120 1277.580 ;
  LAYER metal3 ;
  RECT 0.000 1274.340 1.120 1277.580 ;
  LAYER metal2 ;
  RECT 0.000 1274.340 1.120 1277.580 ;
  LAYER metal1 ;
  RECT 0.000 1274.340 1.120 1277.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1266.500 1.120 1269.740 ;
  LAYER metal3 ;
  RECT 0.000 1266.500 1.120 1269.740 ;
  LAYER metal2 ;
  RECT 0.000 1266.500 1.120 1269.740 ;
  LAYER metal1 ;
  RECT 0.000 1266.500 1.120 1269.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1227.300 1.120 1230.540 ;
  LAYER metal3 ;
  RECT 0.000 1227.300 1.120 1230.540 ;
  LAYER metal2 ;
  RECT 0.000 1227.300 1.120 1230.540 ;
  LAYER metal1 ;
  RECT 0.000 1227.300 1.120 1230.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1219.460 1.120 1222.700 ;
  LAYER metal3 ;
  RECT 0.000 1219.460 1.120 1222.700 ;
  LAYER metal2 ;
  RECT 0.000 1219.460 1.120 1222.700 ;
  LAYER metal1 ;
  RECT 0.000 1219.460 1.120 1222.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1211.620 1.120 1214.860 ;
  LAYER metal3 ;
  RECT 0.000 1211.620 1.120 1214.860 ;
  LAYER metal2 ;
  RECT 0.000 1211.620 1.120 1214.860 ;
  LAYER metal1 ;
  RECT 0.000 1211.620 1.120 1214.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1203.780 1.120 1207.020 ;
  LAYER metal3 ;
  RECT 0.000 1203.780 1.120 1207.020 ;
  LAYER metal2 ;
  RECT 0.000 1203.780 1.120 1207.020 ;
  LAYER metal1 ;
  RECT 0.000 1203.780 1.120 1207.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1195.940 1.120 1199.180 ;
  LAYER metal3 ;
  RECT 0.000 1195.940 1.120 1199.180 ;
  LAYER metal2 ;
  RECT 0.000 1195.940 1.120 1199.180 ;
  LAYER metal1 ;
  RECT 0.000 1195.940 1.120 1199.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1188.100 1.120 1191.340 ;
  LAYER metal3 ;
  RECT 0.000 1188.100 1.120 1191.340 ;
  LAYER metal2 ;
  RECT 0.000 1188.100 1.120 1191.340 ;
  LAYER metal1 ;
  RECT 0.000 1188.100 1.120 1191.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1148.900 1.120 1152.140 ;
  LAYER metal3 ;
  RECT 0.000 1148.900 1.120 1152.140 ;
  LAYER metal2 ;
  RECT 0.000 1148.900 1.120 1152.140 ;
  LAYER metal1 ;
  RECT 0.000 1148.900 1.120 1152.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1141.060 1.120 1144.300 ;
  LAYER metal3 ;
  RECT 0.000 1141.060 1.120 1144.300 ;
  LAYER metal2 ;
  RECT 0.000 1141.060 1.120 1144.300 ;
  LAYER metal1 ;
  RECT 0.000 1141.060 1.120 1144.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1133.220 1.120 1136.460 ;
  LAYER metal3 ;
  RECT 0.000 1133.220 1.120 1136.460 ;
  LAYER metal2 ;
  RECT 0.000 1133.220 1.120 1136.460 ;
  LAYER metal1 ;
  RECT 0.000 1133.220 1.120 1136.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1125.380 1.120 1128.620 ;
  LAYER metal3 ;
  RECT 0.000 1125.380 1.120 1128.620 ;
  LAYER metal2 ;
  RECT 0.000 1125.380 1.120 1128.620 ;
  LAYER metal1 ;
  RECT 0.000 1125.380 1.120 1128.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1117.540 1.120 1120.780 ;
  LAYER metal3 ;
  RECT 0.000 1117.540 1.120 1120.780 ;
  LAYER metal2 ;
  RECT 0.000 1117.540 1.120 1120.780 ;
  LAYER metal1 ;
  RECT 0.000 1117.540 1.120 1120.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1109.700 1.120 1112.940 ;
  LAYER metal3 ;
  RECT 0.000 1109.700 1.120 1112.940 ;
  LAYER metal2 ;
  RECT 0.000 1109.700 1.120 1112.940 ;
  LAYER metal1 ;
  RECT 0.000 1109.700 1.120 1112.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1070.500 1.120 1073.740 ;
  LAYER metal3 ;
  RECT 0.000 1070.500 1.120 1073.740 ;
  LAYER metal2 ;
  RECT 0.000 1070.500 1.120 1073.740 ;
  LAYER metal1 ;
  RECT 0.000 1070.500 1.120 1073.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1062.660 1.120 1065.900 ;
  LAYER metal3 ;
  RECT 0.000 1062.660 1.120 1065.900 ;
  LAYER metal2 ;
  RECT 0.000 1062.660 1.120 1065.900 ;
  LAYER metal1 ;
  RECT 0.000 1062.660 1.120 1065.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1054.820 1.120 1058.060 ;
  LAYER metal3 ;
  RECT 0.000 1054.820 1.120 1058.060 ;
  LAYER metal2 ;
  RECT 0.000 1054.820 1.120 1058.060 ;
  LAYER metal1 ;
  RECT 0.000 1054.820 1.120 1058.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1046.980 1.120 1050.220 ;
  LAYER metal3 ;
  RECT 0.000 1046.980 1.120 1050.220 ;
  LAYER metal2 ;
  RECT 0.000 1046.980 1.120 1050.220 ;
  LAYER metal1 ;
  RECT 0.000 1046.980 1.120 1050.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1039.140 1.120 1042.380 ;
  LAYER metal3 ;
  RECT 0.000 1039.140 1.120 1042.380 ;
  LAYER metal2 ;
  RECT 0.000 1039.140 1.120 1042.380 ;
  LAYER metal1 ;
  RECT 0.000 1039.140 1.120 1042.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1031.300 1.120 1034.540 ;
  LAYER metal3 ;
  RECT 0.000 1031.300 1.120 1034.540 ;
  LAYER metal2 ;
  RECT 0.000 1031.300 1.120 1034.540 ;
  LAYER metal1 ;
  RECT 0.000 1031.300 1.120 1034.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 992.100 1.120 995.340 ;
  LAYER metal3 ;
  RECT 0.000 992.100 1.120 995.340 ;
  LAYER metal2 ;
  RECT 0.000 992.100 1.120 995.340 ;
  LAYER metal1 ;
  RECT 0.000 992.100 1.120 995.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 984.260 1.120 987.500 ;
  LAYER metal3 ;
  RECT 0.000 984.260 1.120 987.500 ;
  LAYER metal2 ;
  RECT 0.000 984.260 1.120 987.500 ;
  LAYER metal1 ;
  RECT 0.000 984.260 1.120 987.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 976.420 1.120 979.660 ;
  LAYER metal3 ;
  RECT 0.000 976.420 1.120 979.660 ;
  LAYER metal2 ;
  RECT 0.000 976.420 1.120 979.660 ;
  LAYER metal1 ;
  RECT 0.000 976.420 1.120 979.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 968.580 1.120 971.820 ;
  LAYER metal3 ;
  RECT 0.000 968.580 1.120 971.820 ;
  LAYER metal2 ;
  RECT 0.000 968.580 1.120 971.820 ;
  LAYER metal1 ;
  RECT 0.000 968.580 1.120 971.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 960.740 1.120 963.980 ;
  LAYER metal3 ;
  RECT 0.000 960.740 1.120 963.980 ;
  LAYER metal2 ;
  RECT 0.000 960.740 1.120 963.980 ;
  LAYER metal1 ;
  RECT 0.000 960.740 1.120 963.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 952.900 1.120 956.140 ;
  LAYER metal3 ;
  RECT 0.000 952.900 1.120 956.140 ;
  LAYER metal2 ;
  RECT 0.000 952.900 1.120 956.140 ;
  LAYER metal1 ;
  RECT 0.000 952.900 1.120 956.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 913.700 1.120 916.940 ;
  LAYER metal3 ;
  RECT 0.000 913.700 1.120 916.940 ;
  LAYER metal2 ;
  RECT 0.000 913.700 1.120 916.940 ;
  LAYER metal1 ;
  RECT 0.000 913.700 1.120 916.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 905.860 1.120 909.100 ;
  LAYER metal3 ;
  RECT 0.000 905.860 1.120 909.100 ;
  LAYER metal2 ;
  RECT 0.000 905.860 1.120 909.100 ;
  LAYER metal1 ;
  RECT 0.000 905.860 1.120 909.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 898.020 1.120 901.260 ;
  LAYER metal3 ;
  RECT 0.000 898.020 1.120 901.260 ;
  LAYER metal2 ;
  RECT 0.000 898.020 1.120 901.260 ;
  LAYER metal1 ;
  RECT 0.000 898.020 1.120 901.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 890.180 1.120 893.420 ;
  LAYER metal3 ;
  RECT 0.000 890.180 1.120 893.420 ;
  LAYER metal2 ;
  RECT 0.000 890.180 1.120 893.420 ;
  LAYER metal1 ;
  RECT 0.000 890.180 1.120 893.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 882.340 1.120 885.580 ;
  LAYER metal3 ;
  RECT 0.000 882.340 1.120 885.580 ;
  LAYER metal2 ;
  RECT 0.000 882.340 1.120 885.580 ;
  LAYER metal1 ;
  RECT 0.000 882.340 1.120 885.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 874.500 1.120 877.740 ;
  LAYER metal3 ;
  RECT 0.000 874.500 1.120 877.740 ;
  LAYER metal2 ;
  RECT 0.000 874.500 1.120 877.740 ;
  LAYER metal1 ;
  RECT 0.000 874.500 1.120 877.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 835.300 1.120 838.540 ;
  LAYER metal3 ;
  RECT 0.000 835.300 1.120 838.540 ;
  LAYER metal2 ;
  RECT 0.000 835.300 1.120 838.540 ;
  LAYER metal1 ;
  RECT 0.000 835.300 1.120 838.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 827.460 1.120 830.700 ;
  LAYER metal3 ;
  RECT 0.000 827.460 1.120 830.700 ;
  LAYER metal2 ;
  RECT 0.000 827.460 1.120 830.700 ;
  LAYER metal1 ;
  RECT 0.000 827.460 1.120 830.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 819.620 1.120 822.860 ;
  LAYER metal3 ;
  RECT 0.000 819.620 1.120 822.860 ;
  LAYER metal2 ;
  RECT 0.000 819.620 1.120 822.860 ;
  LAYER metal1 ;
  RECT 0.000 819.620 1.120 822.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 811.780 1.120 815.020 ;
  LAYER metal3 ;
  RECT 0.000 811.780 1.120 815.020 ;
  LAYER metal2 ;
  RECT 0.000 811.780 1.120 815.020 ;
  LAYER metal1 ;
  RECT 0.000 811.780 1.120 815.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 803.940 1.120 807.180 ;
  LAYER metal3 ;
  RECT 0.000 803.940 1.120 807.180 ;
  LAYER metal2 ;
  RECT 0.000 803.940 1.120 807.180 ;
  LAYER metal1 ;
  RECT 0.000 803.940 1.120 807.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 796.100 1.120 799.340 ;
  LAYER metal3 ;
  RECT 0.000 796.100 1.120 799.340 ;
  LAYER metal2 ;
  RECT 0.000 796.100 1.120 799.340 ;
  LAYER metal1 ;
  RECT 0.000 796.100 1.120 799.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 756.900 1.120 760.140 ;
  LAYER metal3 ;
  RECT 0.000 756.900 1.120 760.140 ;
  LAYER metal2 ;
  RECT 0.000 756.900 1.120 760.140 ;
  LAYER metal1 ;
  RECT 0.000 756.900 1.120 760.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 749.060 1.120 752.300 ;
  LAYER metal3 ;
  RECT 0.000 749.060 1.120 752.300 ;
  LAYER metal2 ;
  RECT 0.000 749.060 1.120 752.300 ;
  LAYER metal1 ;
  RECT 0.000 749.060 1.120 752.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 741.220 1.120 744.460 ;
  LAYER metal3 ;
  RECT 0.000 741.220 1.120 744.460 ;
  LAYER metal2 ;
  RECT 0.000 741.220 1.120 744.460 ;
  LAYER metal1 ;
  RECT 0.000 741.220 1.120 744.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 733.380 1.120 736.620 ;
  LAYER metal3 ;
  RECT 0.000 733.380 1.120 736.620 ;
  LAYER metal2 ;
  RECT 0.000 733.380 1.120 736.620 ;
  LAYER metal1 ;
  RECT 0.000 733.380 1.120 736.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 725.540 1.120 728.780 ;
  LAYER metal3 ;
  RECT 0.000 725.540 1.120 728.780 ;
  LAYER metal2 ;
  RECT 0.000 725.540 1.120 728.780 ;
  LAYER metal1 ;
  RECT 0.000 725.540 1.120 728.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 717.700 1.120 720.940 ;
  LAYER metal3 ;
  RECT 0.000 717.700 1.120 720.940 ;
  LAYER metal2 ;
  RECT 0.000 717.700 1.120 720.940 ;
  LAYER metal1 ;
  RECT 0.000 717.700 1.120 720.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 678.500 1.120 681.740 ;
  LAYER metal3 ;
  RECT 0.000 678.500 1.120 681.740 ;
  LAYER metal2 ;
  RECT 0.000 678.500 1.120 681.740 ;
  LAYER metal1 ;
  RECT 0.000 678.500 1.120 681.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 670.660 1.120 673.900 ;
  LAYER metal3 ;
  RECT 0.000 670.660 1.120 673.900 ;
  LAYER metal2 ;
  RECT 0.000 670.660 1.120 673.900 ;
  LAYER metal1 ;
  RECT 0.000 670.660 1.120 673.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 662.820 1.120 666.060 ;
  LAYER metal3 ;
  RECT 0.000 662.820 1.120 666.060 ;
  LAYER metal2 ;
  RECT 0.000 662.820 1.120 666.060 ;
  LAYER metal1 ;
  RECT 0.000 662.820 1.120 666.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 654.980 1.120 658.220 ;
  LAYER metal3 ;
  RECT 0.000 654.980 1.120 658.220 ;
  LAYER metal2 ;
  RECT 0.000 654.980 1.120 658.220 ;
  LAYER metal1 ;
  RECT 0.000 654.980 1.120 658.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 647.140 1.120 650.380 ;
  LAYER metal3 ;
  RECT 0.000 647.140 1.120 650.380 ;
  LAYER metal2 ;
  RECT 0.000 647.140 1.120 650.380 ;
  LAYER metal1 ;
  RECT 0.000 647.140 1.120 650.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 639.300 1.120 642.540 ;
  LAYER metal3 ;
  RECT 0.000 639.300 1.120 642.540 ;
  LAYER metal2 ;
  RECT 0.000 639.300 1.120 642.540 ;
  LAYER metal1 ;
  RECT 0.000 639.300 1.120 642.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 600.100 1.120 603.340 ;
  LAYER metal3 ;
  RECT 0.000 600.100 1.120 603.340 ;
  LAYER metal2 ;
  RECT 0.000 600.100 1.120 603.340 ;
  LAYER metal1 ;
  RECT 0.000 600.100 1.120 603.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 592.260 1.120 595.500 ;
  LAYER metal3 ;
  RECT 0.000 592.260 1.120 595.500 ;
  LAYER metal2 ;
  RECT 0.000 592.260 1.120 595.500 ;
  LAYER metal1 ;
  RECT 0.000 592.260 1.120 595.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 584.420 1.120 587.660 ;
  LAYER metal3 ;
  RECT 0.000 584.420 1.120 587.660 ;
  LAYER metal2 ;
  RECT 0.000 584.420 1.120 587.660 ;
  LAYER metal1 ;
  RECT 0.000 584.420 1.120 587.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 576.580 1.120 579.820 ;
  LAYER metal3 ;
  RECT 0.000 576.580 1.120 579.820 ;
  LAYER metal2 ;
  RECT 0.000 576.580 1.120 579.820 ;
  LAYER metal1 ;
  RECT 0.000 576.580 1.120 579.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 568.740 1.120 571.980 ;
  LAYER metal3 ;
  RECT 0.000 568.740 1.120 571.980 ;
  LAYER metal2 ;
  RECT 0.000 568.740 1.120 571.980 ;
  LAYER metal1 ;
  RECT 0.000 568.740 1.120 571.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 560.900 1.120 564.140 ;
  LAYER metal3 ;
  RECT 0.000 560.900 1.120 564.140 ;
  LAYER metal2 ;
  RECT 0.000 560.900 1.120 564.140 ;
  LAYER metal1 ;
  RECT 0.000 560.900 1.120 564.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER metal3 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER metal2 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER metal1 ;
  RECT 0.000 521.700 1.120 524.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER metal3 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER metal2 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER metal1 ;
  RECT 0.000 513.860 1.120 517.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER metal3 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER metal2 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER metal1 ;
  RECT 0.000 506.020 1.120 509.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER metal3 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER metal2 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER metal1 ;
  RECT 0.000 498.180 1.120 501.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER metal3 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER metal2 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER metal1 ;
  RECT 0.000 490.340 1.120 493.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER metal3 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER metal2 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER metal1 ;
  RECT 0.000 482.500 1.120 485.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER metal3 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER metal2 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER metal1 ;
  RECT 0.000 443.300 1.120 446.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER metal3 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER metal2 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER metal1 ;
  RECT 0.000 435.460 1.120 438.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER metal3 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER metal2 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER metal1 ;
  RECT 0.000 427.620 1.120 430.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER metal3 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER metal2 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER metal1 ;
  RECT 0.000 419.780 1.120 423.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER metal3 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER metal2 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER metal1 ;
  RECT 0.000 411.940 1.120 415.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER metal3 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER metal2 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER metal1 ;
  RECT 0.000 404.100 1.120 407.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER metal3 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER metal2 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER metal1 ;
  RECT 0.000 364.900 1.120 368.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER metal3 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER metal2 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER metal1 ;
  RECT 0.000 357.060 1.120 360.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER metal3 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER metal2 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER metal1 ;
  RECT 0.000 349.220 1.120 352.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER metal3 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER metal2 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER metal1 ;
  RECT 0.000 341.380 1.120 344.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER metal3 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER metal2 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER metal1 ;
  RECT 0.000 333.540 1.120 336.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER metal3 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER metal2 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER metal1 ;
  RECT 0.000 325.700 1.120 328.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER metal3 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER metal2 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER metal1 ;
  RECT 0.000 286.500 1.120 289.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal3 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal2 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal1 ;
  RECT 0.000 278.660 1.120 281.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal3 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal2 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal1 ;
  RECT 0.000 270.820 1.120 274.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal3 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal2 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal1 ;
  RECT 0.000 262.980 1.120 266.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal3 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal2 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal1 ;
  RECT 0.000 255.140 1.120 258.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal3 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal2 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal1 ;
  RECT 0.000 247.300 1.120 250.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal3 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal2 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal1 ;
  RECT 0.000 208.100 1.120 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1878.380 1390.480 1881.920 1391.600 ;
  LAYER metal3 ;
  RECT 1878.380 1390.480 1881.920 1391.600 ;
  LAYER metal2 ;
  RECT 1878.380 1390.480 1881.920 1391.600 ;
  LAYER metal1 ;
  RECT 1878.380 1390.480 1881.920 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1869.700 1390.480 1873.240 1391.600 ;
  LAYER metal3 ;
  RECT 1869.700 1390.480 1873.240 1391.600 ;
  LAYER metal2 ;
  RECT 1869.700 1390.480 1873.240 1391.600 ;
  LAYER metal1 ;
  RECT 1869.700 1390.480 1873.240 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1861.020 1390.480 1864.560 1391.600 ;
  LAYER metal3 ;
  RECT 1861.020 1390.480 1864.560 1391.600 ;
  LAYER metal2 ;
  RECT 1861.020 1390.480 1864.560 1391.600 ;
  LAYER metal1 ;
  RECT 1861.020 1390.480 1864.560 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1852.340 1390.480 1855.880 1391.600 ;
  LAYER metal3 ;
  RECT 1852.340 1390.480 1855.880 1391.600 ;
  LAYER metal2 ;
  RECT 1852.340 1390.480 1855.880 1391.600 ;
  LAYER metal1 ;
  RECT 1852.340 1390.480 1855.880 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1843.660 1390.480 1847.200 1391.600 ;
  LAYER metal3 ;
  RECT 1843.660 1390.480 1847.200 1391.600 ;
  LAYER metal2 ;
  RECT 1843.660 1390.480 1847.200 1391.600 ;
  LAYER metal1 ;
  RECT 1843.660 1390.480 1847.200 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1834.980 1390.480 1838.520 1391.600 ;
  LAYER metal3 ;
  RECT 1834.980 1390.480 1838.520 1391.600 ;
  LAYER metal2 ;
  RECT 1834.980 1390.480 1838.520 1391.600 ;
  LAYER metal1 ;
  RECT 1834.980 1390.480 1838.520 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1791.580 1390.480 1795.120 1391.600 ;
  LAYER metal3 ;
  RECT 1791.580 1390.480 1795.120 1391.600 ;
  LAYER metal2 ;
  RECT 1791.580 1390.480 1795.120 1391.600 ;
  LAYER metal1 ;
  RECT 1791.580 1390.480 1795.120 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1782.900 1390.480 1786.440 1391.600 ;
  LAYER metal3 ;
  RECT 1782.900 1390.480 1786.440 1391.600 ;
  LAYER metal2 ;
  RECT 1782.900 1390.480 1786.440 1391.600 ;
  LAYER metal1 ;
  RECT 1782.900 1390.480 1786.440 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1774.220 1390.480 1777.760 1391.600 ;
  LAYER metal3 ;
  RECT 1774.220 1390.480 1777.760 1391.600 ;
  LAYER metal2 ;
  RECT 1774.220 1390.480 1777.760 1391.600 ;
  LAYER metal1 ;
  RECT 1774.220 1390.480 1777.760 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1765.540 1390.480 1769.080 1391.600 ;
  LAYER metal3 ;
  RECT 1765.540 1390.480 1769.080 1391.600 ;
  LAYER metal2 ;
  RECT 1765.540 1390.480 1769.080 1391.600 ;
  LAYER metal1 ;
  RECT 1765.540 1390.480 1769.080 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1756.860 1390.480 1760.400 1391.600 ;
  LAYER metal3 ;
  RECT 1756.860 1390.480 1760.400 1391.600 ;
  LAYER metal2 ;
  RECT 1756.860 1390.480 1760.400 1391.600 ;
  LAYER metal1 ;
  RECT 1756.860 1390.480 1760.400 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1748.180 1390.480 1751.720 1391.600 ;
  LAYER metal3 ;
  RECT 1748.180 1390.480 1751.720 1391.600 ;
  LAYER metal2 ;
  RECT 1748.180 1390.480 1751.720 1391.600 ;
  LAYER metal1 ;
  RECT 1748.180 1390.480 1751.720 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1704.780 1390.480 1708.320 1391.600 ;
  LAYER metal3 ;
  RECT 1704.780 1390.480 1708.320 1391.600 ;
  LAYER metal2 ;
  RECT 1704.780 1390.480 1708.320 1391.600 ;
  LAYER metal1 ;
  RECT 1704.780 1390.480 1708.320 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1696.100 1390.480 1699.640 1391.600 ;
  LAYER metal3 ;
  RECT 1696.100 1390.480 1699.640 1391.600 ;
  LAYER metal2 ;
  RECT 1696.100 1390.480 1699.640 1391.600 ;
  LAYER metal1 ;
  RECT 1696.100 1390.480 1699.640 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1687.420 1390.480 1690.960 1391.600 ;
  LAYER metal3 ;
  RECT 1687.420 1390.480 1690.960 1391.600 ;
  LAYER metal2 ;
  RECT 1687.420 1390.480 1690.960 1391.600 ;
  LAYER metal1 ;
  RECT 1687.420 1390.480 1690.960 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1678.740 1390.480 1682.280 1391.600 ;
  LAYER metal3 ;
  RECT 1678.740 1390.480 1682.280 1391.600 ;
  LAYER metal2 ;
  RECT 1678.740 1390.480 1682.280 1391.600 ;
  LAYER metal1 ;
  RECT 1678.740 1390.480 1682.280 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1670.060 1390.480 1673.600 1391.600 ;
  LAYER metal3 ;
  RECT 1670.060 1390.480 1673.600 1391.600 ;
  LAYER metal2 ;
  RECT 1670.060 1390.480 1673.600 1391.600 ;
  LAYER metal1 ;
  RECT 1670.060 1390.480 1673.600 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1661.380 1390.480 1664.920 1391.600 ;
  LAYER metal3 ;
  RECT 1661.380 1390.480 1664.920 1391.600 ;
  LAYER metal2 ;
  RECT 1661.380 1390.480 1664.920 1391.600 ;
  LAYER metal1 ;
  RECT 1661.380 1390.480 1664.920 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1617.980 1390.480 1621.520 1391.600 ;
  LAYER metal3 ;
  RECT 1617.980 1390.480 1621.520 1391.600 ;
  LAYER metal2 ;
  RECT 1617.980 1390.480 1621.520 1391.600 ;
  LAYER metal1 ;
  RECT 1617.980 1390.480 1621.520 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1609.300 1390.480 1612.840 1391.600 ;
  LAYER metal3 ;
  RECT 1609.300 1390.480 1612.840 1391.600 ;
  LAYER metal2 ;
  RECT 1609.300 1390.480 1612.840 1391.600 ;
  LAYER metal1 ;
  RECT 1609.300 1390.480 1612.840 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1600.620 1390.480 1604.160 1391.600 ;
  LAYER metal3 ;
  RECT 1600.620 1390.480 1604.160 1391.600 ;
  LAYER metal2 ;
  RECT 1600.620 1390.480 1604.160 1391.600 ;
  LAYER metal1 ;
  RECT 1600.620 1390.480 1604.160 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1591.940 1390.480 1595.480 1391.600 ;
  LAYER metal3 ;
  RECT 1591.940 1390.480 1595.480 1391.600 ;
  LAYER metal2 ;
  RECT 1591.940 1390.480 1595.480 1391.600 ;
  LAYER metal1 ;
  RECT 1591.940 1390.480 1595.480 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1583.260 1390.480 1586.800 1391.600 ;
  LAYER metal3 ;
  RECT 1583.260 1390.480 1586.800 1391.600 ;
  LAYER metal2 ;
  RECT 1583.260 1390.480 1586.800 1391.600 ;
  LAYER metal1 ;
  RECT 1583.260 1390.480 1586.800 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1574.580 1390.480 1578.120 1391.600 ;
  LAYER metal3 ;
  RECT 1574.580 1390.480 1578.120 1391.600 ;
  LAYER metal2 ;
  RECT 1574.580 1390.480 1578.120 1391.600 ;
  LAYER metal1 ;
  RECT 1574.580 1390.480 1578.120 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1531.180 1390.480 1534.720 1391.600 ;
  LAYER metal3 ;
  RECT 1531.180 1390.480 1534.720 1391.600 ;
  LAYER metal2 ;
  RECT 1531.180 1390.480 1534.720 1391.600 ;
  LAYER metal1 ;
  RECT 1531.180 1390.480 1534.720 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1522.500 1390.480 1526.040 1391.600 ;
  LAYER metal3 ;
  RECT 1522.500 1390.480 1526.040 1391.600 ;
  LAYER metal2 ;
  RECT 1522.500 1390.480 1526.040 1391.600 ;
  LAYER metal1 ;
  RECT 1522.500 1390.480 1526.040 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1513.820 1390.480 1517.360 1391.600 ;
  LAYER metal3 ;
  RECT 1513.820 1390.480 1517.360 1391.600 ;
  LAYER metal2 ;
  RECT 1513.820 1390.480 1517.360 1391.600 ;
  LAYER metal1 ;
  RECT 1513.820 1390.480 1517.360 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1505.140 1390.480 1508.680 1391.600 ;
  LAYER metal3 ;
  RECT 1505.140 1390.480 1508.680 1391.600 ;
  LAYER metal2 ;
  RECT 1505.140 1390.480 1508.680 1391.600 ;
  LAYER metal1 ;
  RECT 1505.140 1390.480 1508.680 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1496.460 1390.480 1500.000 1391.600 ;
  LAYER metal3 ;
  RECT 1496.460 1390.480 1500.000 1391.600 ;
  LAYER metal2 ;
  RECT 1496.460 1390.480 1500.000 1391.600 ;
  LAYER metal1 ;
  RECT 1496.460 1390.480 1500.000 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1487.780 1390.480 1491.320 1391.600 ;
  LAYER metal3 ;
  RECT 1487.780 1390.480 1491.320 1391.600 ;
  LAYER metal2 ;
  RECT 1487.780 1390.480 1491.320 1391.600 ;
  LAYER metal1 ;
  RECT 1487.780 1390.480 1491.320 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1444.380 1390.480 1447.920 1391.600 ;
  LAYER metal3 ;
  RECT 1444.380 1390.480 1447.920 1391.600 ;
  LAYER metal2 ;
  RECT 1444.380 1390.480 1447.920 1391.600 ;
  LAYER metal1 ;
  RECT 1444.380 1390.480 1447.920 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1435.700 1390.480 1439.240 1391.600 ;
  LAYER metal3 ;
  RECT 1435.700 1390.480 1439.240 1391.600 ;
  LAYER metal2 ;
  RECT 1435.700 1390.480 1439.240 1391.600 ;
  LAYER metal1 ;
  RECT 1435.700 1390.480 1439.240 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1427.020 1390.480 1430.560 1391.600 ;
  LAYER metal3 ;
  RECT 1427.020 1390.480 1430.560 1391.600 ;
  LAYER metal2 ;
  RECT 1427.020 1390.480 1430.560 1391.600 ;
  LAYER metal1 ;
  RECT 1427.020 1390.480 1430.560 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1418.340 1390.480 1421.880 1391.600 ;
  LAYER metal3 ;
  RECT 1418.340 1390.480 1421.880 1391.600 ;
  LAYER metal2 ;
  RECT 1418.340 1390.480 1421.880 1391.600 ;
  LAYER metal1 ;
  RECT 1418.340 1390.480 1421.880 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1409.660 1390.480 1413.200 1391.600 ;
  LAYER metal3 ;
  RECT 1409.660 1390.480 1413.200 1391.600 ;
  LAYER metal2 ;
  RECT 1409.660 1390.480 1413.200 1391.600 ;
  LAYER metal1 ;
  RECT 1409.660 1390.480 1413.200 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1400.980 1390.480 1404.520 1391.600 ;
  LAYER metal3 ;
  RECT 1400.980 1390.480 1404.520 1391.600 ;
  LAYER metal2 ;
  RECT 1400.980 1390.480 1404.520 1391.600 ;
  LAYER metal1 ;
  RECT 1400.980 1390.480 1404.520 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1357.580 1390.480 1361.120 1391.600 ;
  LAYER metal3 ;
  RECT 1357.580 1390.480 1361.120 1391.600 ;
  LAYER metal2 ;
  RECT 1357.580 1390.480 1361.120 1391.600 ;
  LAYER metal1 ;
  RECT 1357.580 1390.480 1361.120 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1348.900 1390.480 1352.440 1391.600 ;
  LAYER metal3 ;
  RECT 1348.900 1390.480 1352.440 1391.600 ;
  LAYER metal2 ;
  RECT 1348.900 1390.480 1352.440 1391.600 ;
  LAYER metal1 ;
  RECT 1348.900 1390.480 1352.440 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1340.220 1390.480 1343.760 1391.600 ;
  LAYER metal3 ;
  RECT 1340.220 1390.480 1343.760 1391.600 ;
  LAYER metal2 ;
  RECT 1340.220 1390.480 1343.760 1391.600 ;
  LAYER metal1 ;
  RECT 1340.220 1390.480 1343.760 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1331.540 1390.480 1335.080 1391.600 ;
  LAYER metal3 ;
  RECT 1331.540 1390.480 1335.080 1391.600 ;
  LAYER metal2 ;
  RECT 1331.540 1390.480 1335.080 1391.600 ;
  LAYER metal1 ;
  RECT 1331.540 1390.480 1335.080 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1322.860 1390.480 1326.400 1391.600 ;
  LAYER metal3 ;
  RECT 1322.860 1390.480 1326.400 1391.600 ;
  LAYER metal2 ;
  RECT 1322.860 1390.480 1326.400 1391.600 ;
  LAYER metal1 ;
  RECT 1322.860 1390.480 1326.400 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1314.180 1390.480 1317.720 1391.600 ;
  LAYER metal3 ;
  RECT 1314.180 1390.480 1317.720 1391.600 ;
  LAYER metal2 ;
  RECT 1314.180 1390.480 1317.720 1391.600 ;
  LAYER metal1 ;
  RECT 1314.180 1390.480 1317.720 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1270.780 1390.480 1274.320 1391.600 ;
  LAYER metal3 ;
  RECT 1270.780 1390.480 1274.320 1391.600 ;
  LAYER metal2 ;
  RECT 1270.780 1390.480 1274.320 1391.600 ;
  LAYER metal1 ;
  RECT 1270.780 1390.480 1274.320 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1262.100 1390.480 1265.640 1391.600 ;
  LAYER metal3 ;
  RECT 1262.100 1390.480 1265.640 1391.600 ;
  LAYER metal2 ;
  RECT 1262.100 1390.480 1265.640 1391.600 ;
  LAYER metal1 ;
  RECT 1262.100 1390.480 1265.640 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1253.420 1390.480 1256.960 1391.600 ;
  LAYER metal3 ;
  RECT 1253.420 1390.480 1256.960 1391.600 ;
  LAYER metal2 ;
  RECT 1253.420 1390.480 1256.960 1391.600 ;
  LAYER metal1 ;
  RECT 1253.420 1390.480 1256.960 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1244.740 1390.480 1248.280 1391.600 ;
  LAYER metal3 ;
  RECT 1244.740 1390.480 1248.280 1391.600 ;
  LAYER metal2 ;
  RECT 1244.740 1390.480 1248.280 1391.600 ;
  LAYER metal1 ;
  RECT 1244.740 1390.480 1248.280 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1236.060 1390.480 1239.600 1391.600 ;
  LAYER metal3 ;
  RECT 1236.060 1390.480 1239.600 1391.600 ;
  LAYER metal2 ;
  RECT 1236.060 1390.480 1239.600 1391.600 ;
  LAYER metal1 ;
  RECT 1236.060 1390.480 1239.600 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1227.380 1390.480 1230.920 1391.600 ;
  LAYER metal3 ;
  RECT 1227.380 1390.480 1230.920 1391.600 ;
  LAYER metal2 ;
  RECT 1227.380 1390.480 1230.920 1391.600 ;
  LAYER metal1 ;
  RECT 1227.380 1390.480 1230.920 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1183.980 1390.480 1187.520 1391.600 ;
  LAYER metal3 ;
  RECT 1183.980 1390.480 1187.520 1391.600 ;
  LAYER metal2 ;
  RECT 1183.980 1390.480 1187.520 1391.600 ;
  LAYER metal1 ;
  RECT 1183.980 1390.480 1187.520 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1175.300 1390.480 1178.840 1391.600 ;
  LAYER metal3 ;
  RECT 1175.300 1390.480 1178.840 1391.600 ;
  LAYER metal2 ;
  RECT 1175.300 1390.480 1178.840 1391.600 ;
  LAYER metal1 ;
  RECT 1175.300 1390.480 1178.840 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1166.620 1390.480 1170.160 1391.600 ;
  LAYER metal3 ;
  RECT 1166.620 1390.480 1170.160 1391.600 ;
  LAYER metal2 ;
  RECT 1166.620 1390.480 1170.160 1391.600 ;
  LAYER metal1 ;
  RECT 1166.620 1390.480 1170.160 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1157.940 1390.480 1161.480 1391.600 ;
  LAYER metal3 ;
  RECT 1157.940 1390.480 1161.480 1391.600 ;
  LAYER metal2 ;
  RECT 1157.940 1390.480 1161.480 1391.600 ;
  LAYER metal1 ;
  RECT 1157.940 1390.480 1161.480 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1149.260 1390.480 1152.800 1391.600 ;
  LAYER metal3 ;
  RECT 1149.260 1390.480 1152.800 1391.600 ;
  LAYER metal2 ;
  RECT 1149.260 1390.480 1152.800 1391.600 ;
  LAYER metal1 ;
  RECT 1149.260 1390.480 1152.800 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1140.580 1390.480 1144.120 1391.600 ;
  LAYER metal3 ;
  RECT 1140.580 1390.480 1144.120 1391.600 ;
  LAYER metal2 ;
  RECT 1140.580 1390.480 1144.120 1391.600 ;
  LAYER metal1 ;
  RECT 1140.580 1390.480 1144.120 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1097.180 1390.480 1100.720 1391.600 ;
  LAYER metal3 ;
  RECT 1097.180 1390.480 1100.720 1391.600 ;
  LAYER metal2 ;
  RECT 1097.180 1390.480 1100.720 1391.600 ;
  LAYER metal1 ;
  RECT 1097.180 1390.480 1100.720 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1088.500 1390.480 1092.040 1391.600 ;
  LAYER metal3 ;
  RECT 1088.500 1390.480 1092.040 1391.600 ;
  LAYER metal2 ;
  RECT 1088.500 1390.480 1092.040 1391.600 ;
  LAYER metal1 ;
  RECT 1088.500 1390.480 1092.040 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1079.820 1390.480 1083.360 1391.600 ;
  LAYER metal3 ;
  RECT 1079.820 1390.480 1083.360 1391.600 ;
  LAYER metal2 ;
  RECT 1079.820 1390.480 1083.360 1391.600 ;
  LAYER metal1 ;
  RECT 1079.820 1390.480 1083.360 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1071.140 1390.480 1074.680 1391.600 ;
  LAYER metal3 ;
  RECT 1071.140 1390.480 1074.680 1391.600 ;
  LAYER metal2 ;
  RECT 1071.140 1390.480 1074.680 1391.600 ;
  LAYER metal1 ;
  RECT 1071.140 1390.480 1074.680 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1062.460 1390.480 1066.000 1391.600 ;
  LAYER metal3 ;
  RECT 1062.460 1390.480 1066.000 1391.600 ;
  LAYER metal2 ;
  RECT 1062.460 1390.480 1066.000 1391.600 ;
  LAYER metal1 ;
  RECT 1062.460 1390.480 1066.000 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1053.780 1390.480 1057.320 1391.600 ;
  LAYER metal3 ;
  RECT 1053.780 1390.480 1057.320 1391.600 ;
  LAYER metal2 ;
  RECT 1053.780 1390.480 1057.320 1391.600 ;
  LAYER metal1 ;
  RECT 1053.780 1390.480 1057.320 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1010.380 1390.480 1013.920 1391.600 ;
  LAYER metal3 ;
  RECT 1010.380 1390.480 1013.920 1391.600 ;
  LAYER metal2 ;
  RECT 1010.380 1390.480 1013.920 1391.600 ;
  LAYER metal1 ;
  RECT 1010.380 1390.480 1013.920 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1001.700 1390.480 1005.240 1391.600 ;
  LAYER metal3 ;
  RECT 1001.700 1390.480 1005.240 1391.600 ;
  LAYER metal2 ;
  RECT 1001.700 1390.480 1005.240 1391.600 ;
  LAYER metal1 ;
  RECT 1001.700 1390.480 1005.240 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 993.020 1390.480 996.560 1391.600 ;
  LAYER metal3 ;
  RECT 993.020 1390.480 996.560 1391.600 ;
  LAYER metal2 ;
  RECT 993.020 1390.480 996.560 1391.600 ;
  LAYER metal1 ;
  RECT 993.020 1390.480 996.560 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 984.340 1390.480 987.880 1391.600 ;
  LAYER metal3 ;
  RECT 984.340 1390.480 987.880 1391.600 ;
  LAYER metal2 ;
  RECT 984.340 1390.480 987.880 1391.600 ;
  LAYER metal1 ;
  RECT 984.340 1390.480 987.880 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 975.660 1390.480 979.200 1391.600 ;
  LAYER metal3 ;
  RECT 975.660 1390.480 979.200 1391.600 ;
  LAYER metal2 ;
  RECT 975.660 1390.480 979.200 1391.600 ;
  LAYER metal1 ;
  RECT 975.660 1390.480 979.200 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 966.980 1390.480 970.520 1391.600 ;
  LAYER metal3 ;
  RECT 966.980 1390.480 970.520 1391.600 ;
  LAYER metal2 ;
  RECT 966.980 1390.480 970.520 1391.600 ;
  LAYER metal1 ;
  RECT 966.980 1390.480 970.520 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 923.580 1390.480 927.120 1391.600 ;
  LAYER metal3 ;
  RECT 923.580 1390.480 927.120 1391.600 ;
  LAYER metal2 ;
  RECT 923.580 1390.480 927.120 1391.600 ;
  LAYER metal1 ;
  RECT 923.580 1390.480 927.120 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 914.900 1390.480 918.440 1391.600 ;
  LAYER metal3 ;
  RECT 914.900 1390.480 918.440 1391.600 ;
  LAYER metal2 ;
  RECT 914.900 1390.480 918.440 1391.600 ;
  LAYER metal1 ;
  RECT 914.900 1390.480 918.440 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 906.220 1390.480 909.760 1391.600 ;
  LAYER metal3 ;
  RECT 906.220 1390.480 909.760 1391.600 ;
  LAYER metal2 ;
  RECT 906.220 1390.480 909.760 1391.600 ;
  LAYER metal1 ;
  RECT 906.220 1390.480 909.760 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 897.540 1390.480 901.080 1391.600 ;
  LAYER metal3 ;
  RECT 897.540 1390.480 901.080 1391.600 ;
  LAYER metal2 ;
  RECT 897.540 1390.480 901.080 1391.600 ;
  LAYER metal1 ;
  RECT 897.540 1390.480 901.080 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 888.860 1390.480 892.400 1391.600 ;
  LAYER metal3 ;
  RECT 888.860 1390.480 892.400 1391.600 ;
  LAYER metal2 ;
  RECT 888.860 1390.480 892.400 1391.600 ;
  LAYER metal1 ;
  RECT 888.860 1390.480 892.400 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 880.180 1390.480 883.720 1391.600 ;
  LAYER metal3 ;
  RECT 880.180 1390.480 883.720 1391.600 ;
  LAYER metal2 ;
  RECT 880.180 1390.480 883.720 1391.600 ;
  LAYER metal1 ;
  RECT 880.180 1390.480 883.720 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 836.780 1390.480 840.320 1391.600 ;
  LAYER metal3 ;
  RECT 836.780 1390.480 840.320 1391.600 ;
  LAYER metal2 ;
  RECT 836.780 1390.480 840.320 1391.600 ;
  LAYER metal1 ;
  RECT 836.780 1390.480 840.320 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 828.100 1390.480 831.640 1391.600 ;
  LAYER metal3 ;
  RECT 828.100 1390.480 831.640 1391.600 ;
  LAYER metal2 ;
  RECT 828.100 1390.480 831.640 1391.600 ;
  LAYER metal1 ;
  RECT 828.100 1390.480 831.640 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 819.420 1390.480 822.960 1391.600 ;
  LAYER metal3 ;
  RECT 819.420 1390.480 822.960 1391.600 ;
  LAYER metal2 ;
  RECT 819.420 1390.480 822.960 1391.600 ;
  LAYER metal1 ;
  RECT 819.420 1390.480 822.960 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 810.740 1390.480 814.280 1391.600 ;
  LAYER metal3 ;
  RECT 810.740 1390.480 814.280 1391.600 ;
  LAYER metal2 ;
  RECT 810.740 1390.480 814.280 1391.600 ;
  LAYER metal1 ;
  RECT 810.740 1390.480 814.280 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 802.060 1390.480 805.600 1391.600 ;
  LAYER metal3 ;
  RECT 802.060 1390.480 805.600 1391.600 ;
  LAYER metal2 ;
  RECT 802.060 1390.480 805.600 1391.600 ;
  LAYER metal1 ;
  RECT 802.060 1390.480 805.600 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 793.380 1390.480 796.920 1391.600 ;
  LAYER metal3 ;
  RECT 793.380 1390.480 796.920 1391.600 ;
  LAYER metal2 ;
  RECT 793.380 1390.480 796.920 1391.600 ;
  LAYER metal1 ;
  RECT 793.380 1390.480 796.920 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.980 1390.480 753.520 1391.600 ;
  LAYER metal3 ;
  RECT 749.980 1390.480 753.520 1391.600 ;
  LAYER metal2 ;
  RECT 749.980 1390.480 753.520 1391.600 ;
  LAYER metal1 ;
  RECT 749.980 1390.480 753.520 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 741.300 1390.480 744.840 1391.600 ;
  LAYER metal3 ;
  RECT 741.300 1390.480 744.840 1391.600 ;
  LAYER metal2 ;
  RECT 741.300 1390.480 744.840 1391.600 ;
  LAYER metal1 ;
  RECT 741.300 1390.480 744.840 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 732.620 1390.480 736.160 1391.600 ;
  LAYER metal3 ;
  RECT 732.620 1390.480 736.160 1391.600 ;
  LAYER metal2 ;
  RECT 732.620 1390.480 736.160 1391.600 ;
  LAYER metal1 ;
  RECT 732.620 1390.480 736.160 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 723.940 1390.480 727.480 1391.600 ;
  LAYER metal3 ;
  RECT 723.940 1390.480 727.480 1391.600 ;
  LAYER metal2 ;
  RECT 723.940 1390.480 727.480 1391.600 ;
  LAYER metal1 ;
  RECT 723.940 1390.480 727.480 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 715.260 1390.480 718.800 1391.600 ;
  LAYER metal3 ;
  RECT 715.260 1390.480 718.800 1391.600 ;
  LAYER metal2 ;
  RECT 715.260 1390.480 718.800 1391.600 ;
  LAYER metal1 ;
  RECT 715.260 1390.480 718.800 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 706.580 1390.480 710.120 1391.600 ;
  LAYER metal3 ;
  RECT 706.580 1390.480 710.120 1391.600 ;
  LAYER metal2 ;
  RECT 706.580 1390.480 710.120 1391.600 ;
  LAYER metal1 ;
  RECT 706.580 1390.480 710.120 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 663.180 1390.480 666.720 1391.600 ;
  LAYER metal3 ;
  RECT 663.180 1390.480 666.720 1391.600 ;
  LAYER metal2 ;
  RECT 663.180 1390.480 666.720 1391.600 ;
  LAYER metal1 ;
  RECT 663.180 1390.480 666.720 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 654.500 1390.480 658.040 1391.600 ;
  LAYER metal3 ;
  RECT 654.500 1390.480 658.040 1391.600 ;
  LAYER metal2 ;
  RECT 654.500 1390.480 658.040 1391.600 ;
  LAYER metal1 ;
  RECT 654.500 1390.480 658.040 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 645.820 1390.480 649.360 1391.600 ;
  LAYER metal3 ;
  RECT 645.820 1390.480 649.360 1391.600 ;
  LAYER metal2 ;
  RECT 645.820 1390.480 649.360 1391.600 ;
  LAYER metal1 ;
  RECT 645.820 1390.480 649.360 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 637.140 1390.480 640.680 1391.600 ;
  LAYER metal3 ;
  RECT 637.140 1390.480 640.680 1391.600 ;
  LAYER metal2 ;
  RECT 637.140 1390.480 640.680 1391.600 ;
  LAYER metal1 ;
  RECT 637.140 1390.480 640.680 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 628.460 1390.480 632.000 1391.600 ;
  LAYER metal3 ;
  RECT 628.460 1390.480 632.000 1391.600 ;
  LAYER metal2 ;
  RECT 628.460 1390.480 632.000 1391.600 ;
  LAYER metal1 ;
  RECT 628.460 1390.480 632.000 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 619.780 1390.480 623.320 1391.600 ;
  LAYER metal3 ;
  RECT 619.780 1390.480 623.320 1391.600 ;
  LAYER metal2 ;
  RECT 619.780 1390.480 623.320 1391.600 ;
  LAYER metal1 ;
  RECT 619.780 1390.480 623.320 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 576.380 1390.480 579.920 1391.600 ;
  LAYER metal3 ;
  RECT 576.380 1390.480 579.920 1391.600 ;
  LAYER metal2 ;
  RECT 576.380 1390.480 579.920 1391.600 ;
  LAYER metal1 ;
  RECT 576.380 1390.480 579.920 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 567.700 1390.480 571.240 1391.600 ;
  LAYER metal3 ;
  RECT 567.700 1390.480 571.240 1391.600 ;
  LAYER metal2 ;
  RECT 567.700 1390.480 571.240 1391.600 ;
  LAYER metal1 ;
  RECT 567.700 1390.480 571.240 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 559.020 1390.480 562.560 1391.600 ;
  LAYER metal3 ;
  RECT 559.020 1390.480 562.560 1391.600 ;
  LAYER metal2 ;
  RECT 559.020 1390.480 562.560 1391.600 ;
  LAYER metal1 ;
  RECT 559.020 1390.480 562.560 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 550.340 1390.480 553.880 1391.600 ;
  LAYER metal3 ;
  RECT 550.340 1390.480 553.880 1391.600 ;
  LAYER metal2 ;
  RECT 550.340 1390.480 553.880 1391.600 ;
  LAYER metal1 ;
  RECT 550.340 1390.480 553.880 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 541.660 1390.480 545.200 1391.600 ;
  LAYER metal3 ;
  RECT 541.660 1390.480 545.200 1391.600 ;
  LAYER metal2 ;
  RECT 541.660 1390.480 545.200 1391.600 ;
  LAYER metal1 ;
  RECT 541.660 1390.480 545.200 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 532.980 1390.480 536.520 1391.600 ;
  LAYER metal3 ;
  RECT 532.980 1390.480 536.520 1391.600 ;
  LAYER metal2 ;
  RECT 532.980 1390.480 536.520 1391.600 ;
  LAYER metal1 ;
  RECT 532.980 1390.480 536.520 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 489.580 1390.480 493.120 1391.600 ;
  LAYER metal3 ;
  RECT 489.580 1390.480 493.120 1391.600 ;
  LAYER metal2 ;
  RECT 489.580 1390.480 493.120 1391.600 ;
  LAYER metal1 ;
  RECT 489.580 1390.480 493.120 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 480.900 1390.480 484.440 1391.600 ;
  LAYER metal3 ;
  RECT 480.900 1390.480 484.440 1391.600 ;
  LAYER metal2 ;
  RECT 480.900 1390.480 484.440 1391.600 ;
  LAYER metal1 ;
  RECT 480.900 1390.480 484.440 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 472.220 1390.480 475.760 1391.600 ;
  LAYER metal3 ;
  RECT 472.220 1390.480 475.760 1391.600 ;
  LAYER metal2 ;
  RECT 472.220 1390.480 475.760 1391.600 ;
  LAYER metal1 ;
  RECT 472.220 1390.480 475.760 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 463.540 1390.480 467.080 1391.600 ;
  LAYER metal3 ;
  RECT 463.540 1390.480 467.080 1391.600 ;
  LAYER metal2 ;
  RECT 463.540 1390.480 467.080 1391.600 ;
  LAYER metal1 ;
  RECT 463.540 1390.480 467.080 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 454.860 1390.480 458.400 1391.600 ;
  LAYER metal3 ;
  RECT 454.860 1390.480 458.400 1391.600 ;
  LAYER metal2 ;
  RECT 454.860 1390.480 458.400 1391.600 ;
  LAYER metal1 ;
  RECT 454.860 1390.480 458.400 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 446.180 1390.480 449.720 1391.600 ;
  LAYER metal3 ;
  RECT 446.180 1390.480 449.720 1391.600 ;
  LAYER metal2 ;
  RECT 446.180 1390.480 449.720 1391.600 ;
  LAYER metal1 ;
  RECT 446.180 1390.480 449.720 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 402.780 1390.480 406.320 1391.600 ;
  LAYER metal3 ;
  RECT 402.780 1390.480 406.320 1391.600 ;
  LAYER metal2 ;
  RECT 402.780 1390.480 406.320 1391.600 ;
  LAYER metal1 ;
  RECT 402.780 1390.480 406.320 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 394.100 1390.480 397.640 1391.600 ;
  LAYER metal3 ;
  RECT 394.100 1390.480 397.640 1391.600 ;
  LAYER metal2 ;
  RECT 394.100 1390.480 397.640 1391.600 ;
  LAYER metal1 ;
  RECT 394.100 1390.480 397.640 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 385.420 1390.480 388.960 1391.600 ;
  LAYER metal3 ;
  RECT 385.420 1390.480 388.960 1391.600 ;
  LAYER metal2 ;
  RECT 385.420 1390.480 388.960 1391.600 ;
  LAYER metal1 ;
  RECT 385.420 1390.480 388.960 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 376.740 1390.480 380.280 1391.600 ;
  LAYER metal3 ;
  RECT 376.740 1390.480 380.280 1391.600 ;
  LAYER metal2 ;
  RECT 376.740 1390.480 380.280 1391.600 ;
  LAYER metal1 ;
  RECT 376.740 1390.480 380.280 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 368.060 1390.480 371.600 1391.600 ;
  LAYER metal3 ;
  RECT 368.060 1390.480 371.600 1391.600 ;
  LAYER metal2 ;
  RECT 368.060 1390.480 371.600 1391.600 ;
  LAYER metal1 ;
  RECT 368.060 1390.480 371.600 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 359.380 1390.480 362.920 1391.600 ;
  LAYER metal3 ;
  RECT 359.380 1390.480 362.920 1391.600 ;
  LAYER metal2 ;
  RECT 359.380 1390.480 362.920 1391.600 ;
  LAYER metal1 ;
  RECT 359.380 1390.480 362.920 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.980 1390.480 319.520 1391.600 ;
  LAYER metal3 ;
  RECT 315.980 1390.480 319.520 1391.600 ;
  LAYER metal2 ;
  RECT 315.980 1390.480 319.520 1391.600 ;
  LAYER metal1 ;
  RECT 315.980 1390.480 319.520 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 307.300 1390.480 310.840 1391.600 ;
  LAYER metal3 ;
  RECT 307.300 1390.480 310.840 1391.600 ;
  LAYER metal2 ;
  RECT 307.300 1390.480 310.840 1391.600 ;
  LAYER metal1 ;
  RECT 307.300 1390.480 310.840 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 298.620 1390.480 302.160 1391.600 ;
  LAYER metal3 ;
  RECT 298.620 1390.480 302.160 1391.600 ;
  LAYER metal2 ;
  RECT 298.620 1390.480 302.160 1391.600 ;
  LAYER metal1 ;
  RECT 298.620 1390.480 302.160 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 289.940 1390.480 293.480 1391.600 ;
  LAYER metal3 ;
  RECT 289.940 1390.480 293.480 1391.600 ;
  LAYER metal2 ;
  RECT 289.940 1390.480 293.480 1391.600 ;
  LAYER metal1 ;
  RECT 289.940 1390.480 293.480 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 281.260 1390.480 284.800 1391.600 ;
  LAYER metal3 ;
  RECT 281.260 1390.480 284.800 1391.600 ;
  LAYER metal2 ;
  RECT 281.260 1390.480 284.800 1391.600 ;
  LAYER metal1 ;
  RECT 281.260 1390.480 284.800 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 272.580 1390.480 276.120 1391.600 ;
  LAYER metal3 ;
  RECT 272.580 1390.480 276.120 1391.600 ;
  LAYER metal2 ;
  RECT 272.580 1390.480 276.120 1391.600 ;
  LAYER metal1 ;
  RECT 272.580 1390.480 276.120 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.180 1390.480 232.720 1391.600 ;
  LAYER metal3 ;
  RECT 229.180 1390.480 232.720 1391.600 ;
  LAYER metal2 ;
  RECT 229.180 1390.480 232.720 1391.600 ;
  LAYER metal1 ;
  RECT 229.180 1390.480 232.720 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 220.500 1390.480 224.040 1391.600 ;
  LAYER metal3 ;
  RECT 220.500 1390.480 224.040 1391.600 ;
  LAYER metal2 ;
  RECT 220.500 1390.480 224.040 1391.600 ;
  LAYER metal1 ;
  RECT 220.500 1390.480 224.040 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 211.820 1390.480 215.360 1391.600 ;
  LAYER metal3 ;
  RECT 211.820 1390.480 215.360 1391.600 ;
  LAYER metal2 ;
  RECT 211.820 1390.480 215.360 1391.600 ;
  LAYER metal1 ;
  RECT 211.820 1390.480 215.360 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 203.140 1390.480 206.680 1391.600 ;
  LAYER metal3 ;
  RECT 203.140 1390.480 206.680 1391.600 ;
  LAYER metal2 ;
  RECT 203.140 1390.480 206.680 1391.600 ;
  LAYER metal1 ;
  RECT 203.140 1390.480 206.680 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 194.460 1390.480 198.000 1391.600 ;
  LAYER metal3 ;
  RECT 194.460 1390.480 198.000 1391.600 ;
  LAYER metal2 ;
  RECT 194.460 1390.480 198.000 1391.600 ;
  LAYER metal1 ;
  RECT 194.460 1390.480 198.000 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 185.780 1390.480 189.320 1391.600 ;
  LAYER metal3 ;
  RECT 185.780 1390.480 189.320 1391.600 ;
  LAYER metal2 ;
  RECT 185.780 1390.480 189.320 1391.600 ;
  LAYER metal1 ;
  RECT 185.780 1390.480 189.320 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.380 1390.480 145.920 1391.600 ;
  LAYER metal3 ;
  RECT 142.380 1390.480 145.920 1391.600 ;
  LAYER metal2 ;
  RECT 142.380 1390.480 145.920 1391.600 ;
  LAYER metal1 ;
  RECT 142.380 1390.480 145.920 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 133.700 1390.480 137.240 1391.600 ;
  LAYER metal3 ;
  RECT 133.700 1390.480 137.240 1391.600 ;
  LAYER metal2 ;
  RECT 133.700 1390.480 137.240 1391.600 ;
  LAYER metal1 ;
  RECT 133.700 1390.480 137.240 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 125.020 1390.480 128.560 1391.600 ;
  LAYER metal3 ;
  RECT 125.020 1390.480 128.560 1391.600 ;
  LAYER metal2 ;
  RECT 125.020 1390.480 128.560 1391.600 ;
  LAYER metal1 ;
  RECT 125.020 1390.480 128.560 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 116.340 1390.480 119.880 1391.600 ;
  LAYER metal3 ;
  RECT 116.340 1390.480 119.880 1391.600 ;
  LAYER metal2 ;
  RECT 116.340 1390.480 119.880 1391.600 ;
  LAYER metal1 ;
  RECT 116.340 1390.480 119.880 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.660 1390.480 111.200 1391.600 ;
  LAYER metal3 ;
  RECT 107.660 1390.480 111.200 1391.600 ;
  LAYER metal2 ;
  RECT 107.660 1390.480 111.200 1391.600 ;
  LAYER metal1 ;
  RECT 107.660 1390.480 111.200 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 98.980 1390.480 102.520 1391.600 ;
  LAYER metal3 ;
  RECT 98.980 1390.480 102.520 1391.600 ;
  LAYER metal2 ;
  RECT 98.980 1390.480 102.520 1391.600 ;
  LAYER metal1 ;
  RECT 98.980 1390.480 102.520 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 55.580 1390.480 59.120 1391.600 ;
  LAYER metal3 ;
  RECT 55.580 1390.480 59.120 1391.600 ;
  LAYER metal2 ;
  RECT 55.580 1390.480 59.120 1391.600 ;
  LAYER metal1 ;
  RECT 55.580 1390.480 59.120 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 46.900 1390.480 50.440 1391.600 ;
  LAYER metal3 ;
  RECT 46.900 1390.480 50.440 1391.600 ;
  LAYER metal2 ;
  RECT 46.900 1390.480 50.440 1391.600 ;
  LAYER metal1 ;
  RECT 46.900 1390.480 50.440 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 38.220 1390.480 41.760 1391.600 ;
  LAYER metal3 ;
  RECT 38.220 1390.480 41.760 1391.600 ;
  LAYER metal2 ;
  RECT 38.220 1390.480 41.760 1391.600 ;
  LAYER metal1 ;
  RECT 38.220 1390.480 41.760 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 29.540 1390.480 33.080 1391.600 ;
  LAYER metal3 ;
  RECT 29.540 1390.480 33.080 1391.600 ;
  LAYER metal2 ;
  RECT 29.540 1390.480 33.080 1391.600 ;
  LAYER metal1 ;
  RECT 29.540 1390.480 33.080 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 20.860 1390.480 24.400 1391.600 ;
  LAYER metal3 ;
  RECT 20.860 1390.480 24.400 1391.600 ;
  LAYER metal2 ;
  RECT 20.860 1390.480 24.400 1391.600 ;
  LAYER metal1 ;
  RECT 20.860 1390.480 24.400 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.180 1390.480 15.720 1391.600 ;
  LAYER metal3 ;
  RECT 12.180 1390.480 15.720 1391.600 ;
  LAYER metal2 ;
  RECT 12.180 1390.480 15.720 1391.600 ;
  LAYER metal1 ;
  RECT 12.180 1390.480 15.720 1391.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1869.700 0.000 1873.240 1.120 ;
  LAYER metal3 ;
  RECT 1869.700 0.000 1873.240 1.120 ;
  LAYER metal2 ;
  RECT 1869.700 0.000 1873.240 1.120 ;
  LAYER metal1 ;
  RECT 1869.700 0.000 1873.240 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1861.020 0.000 1864.560 1.120 ;
  LAYER metal3 ;
  RECT 1861.020 0.000 1864.560 1.120 ;
  LAYER metal2 ;
  RECT 1861.020 0.000 1864.560 1.120 ;
  LAYER metal1 ;
  RECT 1861.020 0.000 1864.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1852.340 0.000 1855.880 1.120 ;
  LAYER metal3 ;
  RECT 1852.340 0.000 1855.880 1.120 ;
  LAYER metal2 ;
  RECT 1852.340 0.000 1855.880 1.120 ;
  LAYER metal1 ;
  RECT 1852.340 0.000 1855.880 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1843.660 0.000 1847.200 1.120 ;
  LAYER metal3 ;
  RECT 1843.660 0.000 1847.200 1.120 ;
  LAYER metal2 ;
  RECT 1843.660 0.000 1847.200 1.120 ;
  LAYER metal1 ;
  RECT 1843.660 0.000 1847.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1834.980 0.000 1838.520 1.120 ;
  LAYER metal3 ;
  RECT 1834.980 0.000 1838.520 1.120 ;
  LAYER metal2 ;
  RECT 1834.980 0.000 1838.520 1.120 ;
  LAYER metal1 ;
  RECT 1834.980 0.000 1838.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
  LAYER metal3 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
  LAYER metal2 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
  LAYER metal1 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1765.540 0.000 1769.080 1.120 ;
  LAYER metal3 ;
  RECT 1765.540 0.000 1769.080 1.120 ;
  LAYER metal2 ;
  RECT 1765.540 0.000 1769.080 1.120 ;
  LAYER metal1 ;
  RECT 1765.540 0.000 1769.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1756.860 0.000 1760.400 1.120 ;
  LAYER metal3 ;
  RECT 1756.860 0.000 1760.400 1.120 ;
  LAYER metal2 ;
  RECT 1756.860 0.000 1760.400 1.120 ;
  LAYER metal1 ;
  RECT 1756.860 0.000 1760.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1748.180 0.000 1751.720 1.120 ;
  LAYER metal3 ;
  RECT 1748.180 0.000 1751.720 1.120 ;
  LAYER metal2 ;
  RECT 1748.180 0.000 1751.720 1.120 ;
  LAYER metal1 ;
  RECT 1748.180 0.000 1751.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1739.500 0.000 1743.040 1.120 ;
  LAYER metal3 ;
  RECT 1739.500 0.000 1743.040 1.120 ;
  LAYER metal2 ;
  RECT 1739.500 0.000 1743.040 1.120 ;
  LAYER metal1 ;
  RECT 1739.500 0.000 1743.040 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1730.820 0.000 1734.360 1.120 ;
  LAYER metal3 ;
  RECT 1730.820 0.000 1734.360 1.120 ;
  LAYER metal2 ;
  RECT 1730.820 0.000 1734.360 1.120 ;
  LAYER metal1 ;
  RECT 1730.820 0.000 1734.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1722.140 0.000 1725.680 1.120 ;
  LAYER metal3 ;
  RECT 1722.140 0.000 1725.680 1.120 ;
  LAYER metal2 ;
  RECT 1722.140 0.000 1725.680 1.120 ;
  LAYER metal1 ;
  RECT 1722.140 0.000 1725.680 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1661.380 0.000 1664.920 1.120 ;
  LAYER metal3 ;
  RECT 1661.380 0.000 1664.920 1.120 ;
  LAYER metal2 ;
  RECT 1661.380 0.000 1664.920 1.120 ;
  LAYER metal1 ;
  RECT 1661.380 0.000 1664.920 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1652.700 0.000 1656.240 1.120 ;
  LAYER metal3 ;
  RECT 1652.700 0.000 1656.240 1.120 ;
  LAYER metal2 ;
  RECT 1652.700 0.000 1656.240 1.120 ;
  LAYER metal1 ;
  RECT 1652.700 0.000 1656.240 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1644.020 0.000 1647.560 1.120 ;
  LAYER metal3 ;
  RECT 1644.020 0.000 1647.560 1.120 ;
  LAYER metal2 ;
  RECT 1644.020 0.000 1647.560 1.120 ;
  LAYER metal1 ;
  RECT 1644.020 0.000 1647.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1635.340 0.000 1638.880 1.120 ;
  LAYER metal3 ;
  RECT 1635.340 0.000 1638.880 1.120 ;
  LAYER metal2 ;
  RECT 1635.340 0.000 1638.880 1.120 ;
  LAYER metal1 ;
  RECT 1635.340 0.000 1638.880 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1626.660 0.000 1630.200 1.120 ;
  LAYER metal3 ;
  RECT 1626.660 0.000 1630.200 1.120 ;
  LAYER metal2 ;
  RECT 1626.660 0.000 1630.200 1.120 ;
  LAYER metal1 ;
  RECT 1626.660 0.000 1630.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1617.980 0.000 1621.520 1.120 ;
  LAYER metal3 ;
  RECT 1617.980 0.000 1621.520 1.120 ;
  LAYER metal2 ;
  RECT 1617.980 0.000 1621.520 1.120 ;
  LAYER metal1 ;
  RECT 1617.980 0.000 1621.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1556.600 0.000 1560.140 1.120 ;
  LAYER metal3 ;
  RECT 1556.600 0.000 1560.140 1.120 ;
  LAYER metal2 ;
  RECT 1556.600 0.000 1560.140 1.120 ;
  LAYER metal1 ;
  RECT 1556.600 0.000 1560.140 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1547.920 0.000 1551.460 1.120 ;
  LAYER metal3 ;
  RECT 1547.920 0.000 1551.460 1.120 ;
  LAYER metal2 ;
  RECT 1547.920 0.000 1551.460 1.120 ;
  LAYER metal1 ;
  RECT 1547.920 0.000 1551.460 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1539.240 0.000 1542.780 1.120 ;
  LAYER metal3 ;
  RECT 1539.240 0.000 1542.780 1.120 ;
  LAYER metal2 ;
  RECT 1539.240 0.000 1542.780 1.120 ;
  LAYER metal1 ;
  RECT 1539.240 0.000 1542.780 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1530.560 0.000 1534.100 1.120 ;
  LAYER metal3 ;
  RECT 1530.560 0.000 1534.100 1.120 ;
  LAYER metal2 ;
  RECT 1530.560 0.000 1534.100 1.120 ;
  LAYER metal1 ;
  RECT 1530.560 0.000 1534.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1521.880 0.000 1525.420 1.120 ;
  LAYER metal3 ;
  RECT 1521.880 0.000 1525.420 1.120 ;
  LAYER metal2 ;
  RECT 1521.880 0.000 1525.420 1.120 ;
  LAYER metal1 ;
  RECT 1521.880 0.000 1525.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1513.200 0.000 1516.740 1.120 ;
  LAYER metal3 ;
  RECT 1513.200 0.000 1516.740 1.120 ;
  LAYER metal2 ;
  RECT 1513.200 0.000 1516.740 1.120 ;
  LAYER metal1 ;
  RECT 1513.200 0.000 1516.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1452.440 0.000 1455.980 1.120 ;
  LAYER metal3 ;
  RECT 1452.440 0.000 1455.980 1.120 ;
  LAYER metal2 ;
  RECT 1452.440 0.000 1455.980 1.120 ;
  LAYER metal1 ;
  RECT 1452.440 0.000 1455.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1443.760 0.000 1447.300 1.120 ;
  LAYER metal3 ;
  RECT 1443.760 0.000 1447.300 1.120 ;
  LAYER metal2 ;
  RECT 1443.760 0.000 1447.300 1.120 ;
  LAYER metal1 ;
  RECT 1443.760 0.000 1447.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1435.080 0.000 1438.620 1.120 ;
  LAYER metal3 ;
  RECT 1435.080 0.000 1438.620 1.120 ;
  LAYER metal2 ;
  RECT 1435.080 0.000 1438.620 1.120 ;
  LAYER metal1 ;
  RECT 1435.080 0.000 1438.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal3 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal2 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal1 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1417.720 0.000 1421.260 1.120 ;
  LAYER metal3 ;
  RECT 1417.720 0.000 1421.260 1.120 ;
  LAYER metal2 ;
  RECT 1417.720 0.000 1421.260 1.120 ;
  LAYER metal1 ;
  RECT 1417.720 0.000 1421.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1409.040 0.000 1412.580 1.120 ;
  LAYER metal3 ;
  RECT 1409.040 0.000 1412.580 1.120 ;
  LAYER metal2 ;
  RECT 1409.040 0.000 1412.580 1.120 ;
  LAYER metal1 ;
  RECT 1409.040 0.000 1412.580 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1361.920 0.000 1365.460 1.120 ;
  LAYER metal3 ;
  RECT 1361.920 0.000 1365.460 1.120 ;
  LAYER metal2 ;
  RECT 1361.920 0.000 1365.460 1.120 ;
  LAYER metal1 ;
  RECT 1361.920 0.000 1365.460 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1339.600 0.000 1343.140 1.120 ;
  LAYER metal3 ;
  RECT 1339.600 0.000 1343.140 1.120 ;
  LAYER metal2 ;
  RECT 1339.600 0.000 1343.140 1.120 ;
  LAYER metal1 ;
  RECT 1339.600 0.000 1343.140 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1330.920 0.000 1334.460 1.120 ;
  LAYER metal3 ;
  RECT 1330.920 0.000 1334.460 1.120 ;
  LAYER metal2 ;
  RECT 1330.920 0.000 1334.460 1.120 ;
  LAYER metal1 ;
  RECT 1330.920 0.000 1334.460 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1322.240 0.000 1325.780 1.120 ;
  LAYER metal3 ;
  RECT 1322.240 0.000 1325.780 1.120 ;
  LAYER metal2 ;
  RECT 1322.240 0.000 1325.780 1.120 ;
  LAYER metal1 ;
  RECT 1322.240 0.000 1325.780 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1313.560 0.000 1317.100 1.120 ;
  LAYER metal3 ;
  RECT 1313.560 0.000 1317.100 1.120 ;
  LAYER metal2 ;
  RECT 1313.560 0.000 1317.100 1.120 ;
  LAYER metal1 ;
  RECT 1313.560 0.000 1317.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1304.880 0.000 1308.420 1.120 ;
  LAYER metal3 ;
  RECT 1304.880 0.000 1308.420 1.120 ;
  LAYER metal2 ;
  RECT 1304.880 0.000 1308.420 1.120 ;
  LAYER metal1 ;
  RECT 1304.880 0.000 1308.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1261.480 0.000 1265.020 1.120 ;
  LAYER metal3 ;
  RECT 1261.480 0.000 1265.020 1.120 ;
  LAYER metal2 ;
  RECT 1261.480 0.000 1265.020 1.120 ;
  LAYER metal1 ;
  RECT 1261.480 0.000 1265.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1248.460 0.000 1252.000 1.120 ;
  LAYER metal3 ;
  RECT 1248.460 0.000 1252.000 1.120 ;
  LAYER metal2 ;
  RECT 1248.460 0.000 1252.000 1.120 ;
  LAYER metal1 ;
  RECT 1248.460 0.000 1252.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1226.140 0.000 1229.680 1.120 ;
  LAYER metal3 ;
  RECT 1226.140 0.000 1229.680 1.120 ;
  LAYER metal2 ;
  RECT 1226.140 0.000 1229.680 1.120 ;
  LAYER metal1 ;
  RECT 1226.140 0.000 1229.680 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1217.460 0.000 1221.000 1.120 ;
  LAYER metal3 ;
  RECT 1217.460 0.000 1221.000 1.120 ;
  LAYER metal2 ;
  RECT 1217.460 0.000 1221.000 1.120 ;
  LAYER metal1 ;
  RECT 1217.460 0.000 1221.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1208.780 0.000 1212.320 1.120 ;
  LAYER metal3 ;
  RECT 1208.780 0.000 1212.320 1.120 ;
  LAYER metal2 ;
  RECT 1208.780 0.000 1212.320 1.120 ;
  LAYER metal1 ;
  RECT 1208.780 0.000 1212.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1200.100 0.000 1203.640 1.120 ;
  LAYER metal3 ;
  RECT 1200.100 0.000 1203.640 1.120 ;
  LAYER metal2 ;
  RECT 1200.100 0.000 1203.640 1.120 ;
  LAYER metal1 ;
  RECT 1200.100 0.000 1203.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1156.700 0.000 1160.240 1.120 ;
  LAYER metal3 ;
  RECT 1156.700 0.000 1160.240 1.120 ;
  LAYER metal2 ;
  RECT 1156.700 0.000 1160.240 1.120 ;
  LAYER metal1 ;
  RECT 1156.700 0.000 1160.240 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal3 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal2 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal1 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1135.620 0.000 1139.160 1.120 ;
  LAYER metal3 ;
  RECT 1135.620 0.000 1139.160 1.120 ;
  LAYER metal2 ;
  RECT 1135.620 0.000 1139.160 1.120 ;
  LAYER metal1 ;
  RECT 1135.620 0.000 1139.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1113.300 0.000 1116.840 1.120 ;
  LAYER metal3 ;
  RECT 1113.300 0.000 1116.840 1.120 ;
  LAYER metal2 ;
  RECT 1113.300 0.000 1116.840 1.120 ;
  LAYER metal1 ;
  RECT 1113.300 0.000 1116.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1104.620 0.000 1108.160 1.120 ;
  LAYER metal3 ;
  RECT 1104.620 0.000 1108.160 1.120 ;
  LAYER metal2 ;
  RECT 1104.620 0.000 1108.160 1.120 ;
  LAYER metal1 ;
  RECT 1104.620 0.000 1108.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1095.940 0.000 1099.480 1.120 ;
  LAYER metal3 ;
  RECT 1095.940 0.000 1099.480 1.120 ;
  LAYER metal2 ;
  RECT 1095.940 0.000 1099.480 1.120 ;
  LAYER metal1 ;
  RECT 1095.940 0.000 1099.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1052.540 0.000 1056.080 1.120 ;
  LAYER metal3 ;
  RECT 1052.540 0.000 1056.080 1.120 ;
  LAYER metal2 ;
  RECT 1052.540 0.000 1056.080 1.120 ;
  LAYER metal1 ;
  RECT 1052.540 0.000 1056.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1043.860 0.000 1047.400 1.120 ;
  LAYER metal3 ;
  RECT 1043.860 0.000 1047.400 1.120 ;
  LAYER metal2 ;
  RECT 1043.860 0.000 1047.400 1.120 ;
  LAYER metal1 ;
  RECT 1043.860 0.000 1047.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1035.180 0.000 1038.720 1.120 ;
  LAYER metal3 ;
  RECT 1035.180 0.000 1038.720 1.120 ;
  LAYER metal2 ;
  RECT 1035.180 0.000 1038.720 1.120 ;
  LAYER metal1 ;
  RECT 1035.180 0.000 1038.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal3 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal2 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal1 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 986.200 0.000 989.740 1.120 ;
  LAYER metal3 ;
  RECT 986.200 0.000 989.740 1.120 ;
  LAYER metal2 ;
  RECT 986.200 0.000 989.740 1.120 ;
  LAYER metal1 ;
  RECT 986.200 0.000 989.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 973.180 0.000 976.720 1.120 ;
  LAYER metal3 ;
  RECT 973.180 0.000 976.720 1.120 ;
  LAYER metal2 ;
  RECT 973.180 0.000 976.720 1.120 ;
  LAYER metal1 ;
  RECT 973.180 0.000 976.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 891.960 0.000 895.500 1.120 ;
  LAYER metal3 ;
  RECT 891.960 0.000 895.500 1.120 ;
  LAYER metal2 ;
  RECT 891.960 0.000 895.500 1.120 ;
  LAYER metal1 ;
  RECT 891.960 0.000 895.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 883.280 0.000 886.820 1.120 ;
  LAYER metal3 ;
  RECT 883.280 0.000 886.820 1.120 ;
  LAYER metal2 ;
  RECT 883.280 0.000 886.820 1.120 ;
  LAYER metal1 ;
  RECT 883.280 0.000 886.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 874.600 0.000 878.140 1.120 ;
  LAYER metal3 ;
  RECT 874.600 0.000 878.140 1.120 ;
  LAYER metal2 ;
  RECT 874.600 0.000 878.140 1.120 ;
  LAYER metal1 ;
  RECT 874.600 0.000 878.140 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal3 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal2 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal1 ;
  RECT 865.920 0.000 869.460 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 857.240 0.000 860.780 1.120 ;
  LAYER metal3 ;
  RECT 857.240 0.000 860.780 1.120 ;
  LAYER metal2 ;
  RECT 857.240 0.000 860.780 1.120 ;
  LAYER metal1 ;
  RECT 857.240 0.000 860.780 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 848.560 0.000 852.100 1.120 ;
  LAYER metal3 ;
  RECT 848.560 0.000 852.100 1.120 ;
  LAYER metal2 ;
  RECT 848.560 0.000 852.100 1.120 ;
  LAYER metal1 ;
  RECT 848.560 0.000 852.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 787.800 0.000 791.340 1.120 ;
  LAYER metal3 ;
  RECT 787.800 0.000 791.340 1.120 ;
  LAYER metal2 ;
  RECT 787.800 0.000 791.340 1.120 ;
  LAYER metal1 ;
  RECT 787.800 0.000 791.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 779.120 0.000 782.660 1.120 ;
  LAYER metal3 ;
  RECT 779.120 0.000 782.660 1.120 ;
  LAYER metal2 ;
  RECT 779.120 0.000 782.660 1.120 ;
  LAYER metal1 ;
  RECT 779.120 0.000 782.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 770.440 0.000 773.980 1.120 ;
  LAYER metal3 ;
  RECT 770.440 0.000 773.980 1.120 ;
  LAYER metal2 ;
  RECT 770.440 0.000 773.980 1.120 ;
  LAYER metal1 ;
  RECT 770.440 0.000 773.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 761.760 0.000 765.300 1.120 ;
  LAYER metal3 ;
  RECT 761.760 0.000 765.300 1.120 ;
  LAYER metal2 ;
  RECT 761.760 0.000 765.300 1.120 ;
  LAYER metal1 ;
  RECT 761.760 0.000 765.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 753.080 0.000 756.620 1.120 ;
  LAYER metal3 ;
  RECT 753.080 0.000 756.620 1.120 ;
  LAYER metal2 ;
  RECT 753.080 0.000 756.620 1.120 ;
  LAYER metal1 ;
  RECT 753.080 0.000 756.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 744.400 0.000 747.940 1.120 ;
  LAYER metal3 ;
  RECT 744.400 0.000 747.940 1.120 ;
  LAYER metal2 ;
  RECT 744.400 0.000 747.940 1.120 ;
  LAYER metal1 ;
  RECT 744.400 0.000 747.940 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal3 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal2 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal1 ;
  RECT 683.020 0.000 686.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal3 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal2 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal1 ;
  RECT 674.340 0.000 677.880 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal3 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal2 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal1 ;
  RECT 665.660 0.000 669.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal3 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal2 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal1 ;
  RECT 656.980 0.000 660.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 648.300 0.000 651.840 1.120 ;
  LAYER metal3 ;
  RECT 648.300 0.000 651.840 1.120 ;
  LAYER metal2 ;
  RECT 648.300 0.000 651.840 1.120 ;
  LAYER metal1 ;
  RECT 648.300 0.000 651.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 639.620 0.000 643.160 1.120 ;
  LAYER metal3 ;
  RECT 639.620 0.000 643.160 1.120 ;
  LAYER metal2 ;
  RECT 639.620 0.000 643.160 1.120 ;
  LAYER metal1 ;
  RECT 639.620 0.000 643.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 592.500 0.000 596.040 1.120 ;
  LAYER metal3 ;
  RECT 592.500 0.000 596.040 1.120 ;
  LAYER metal2 ;
  RECT 592.500 0.000 596.040 1.120 ;
  LAYER metal1 ;
  RECT 592.500 0.000 596.040 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal3 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal2 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal1 ;
  RECT 570.180 0.000 573.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 561.500 0.000 565.040 1.120 ;
  LAYER metal3 ;
  RECT 561.500 0.000 565.040 1.120 ;
  LAYER metal2 ;
  RECT 561.500 0.000 565.040 1.120 ;
  LAYER metal1 ;
  RECT 561.500 0.000 565.040 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal3 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal2 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal1 ;
  RECT 552.820 0.000 556.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 544.140 0.000 547.680 1.120 ;
  LAYER metal3 ;
  RECT 544.140 0.000 547.680 1.120 ;
  LAYER metal2 ;
  RECT 544.140 0.000 547.680 1.120 ;
  LAYER metal1 ;
  RECT 544.140 0.000 547.680 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 535.460 0.000 539.000 1.120 ;
  LAYER metal3 ;
  RECT 535.460 0.000 539.000 1.120 ;
  LAYER metal2 ;
  RECT 535.460 0.000 539.000 1.120 ;
  LAYER metal1 ;
  RECT 535.460 0.000 539.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 492.060 0.000 495.600 1.120 ;
  LAYER metal3 ;
  RECT 492.060 0.000 495.600 1.120 ;
  LAYER metal2 ;
  RECT 492.060 0.000 495.600 1.120 ;
  LAYER metal1 ;
  RECT 492.060 0.000 495.600 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER metal3 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER metal2 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER metal1 ;
  RECT 479.040 0.000 482.580 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 457.340 0.000 460.880 1.120 ;
  LAYER metal3 ;
  RECT 457.340 0.000 460.880 1.120 ;
  LAYER metal2 ;
  RECT 457.340 0.000 460.880 1.120 ;
  LAYER metal1 ;
  RECT 457.340 0.000 460.880 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 448.660 0.000 452.200 1.120 ;
  LAYER metal3 ;
  RECT 448.660 0.000 452.200 1.120 ;
  LAYER metal2 ;
  RECT 448.660 0.000 452.200 1.120 ;
  LAYER metal1 ;
  RECT 448.660 0.000 452.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER metal3 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER metal2 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER metal1 ;
  RECT 439.980 0.000 443.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal3 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal2 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal1 ;
  RECT 431.300 0.000 434.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 387.900 0.000 391.440 1.120 ;
  LAYER metal3 ;
  RECT 387.900 0.000 391.440 1.120 ;
  LAYER metal2 ;
  RECT 387.900 0.000 391.440 1.120 ;
  LAYER metal1 ;
  RECT 387.900 0.000 391.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 379.220 0.000 382.760 1.120 ;
  LAYER metal3 ;
  RECT 379.220 0.000 382.760 1.120 ;
  LAYER metal2 ;
  RECT 379.220 0.000 382.760 1.120 ;
  LAYER metal1 ;
  RECT 379.220 0.000 382.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER metal3 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER metal2 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER metal1 ;
  RECT 366.200 0.000 369.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 343.880 0.000 347.420 1.120 ;
  LAYER metal3 ;
  RECT 343.880 0.000 347.420 1.120 ;
  LAYER metal2 ;
  RECT 343.880 0.000 347.420 1.120 ;
  LAYER metal1 ;
  RECT 343.880 0.000 347.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 335.200 0.000 338.740 1.120 ;
  LAYER metal3 ;
  RECT 335.200 0.000 338.740 1.120 ;
  LAYER metal2 ;
  RECT 335.200 0.000 338.740 1.120 ;
  LAYER metal1 ;
  RECT 335.200 0.000 338.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal3 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal2 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal1 ;
  RECT 326.520 0.000 330.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal3 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal2 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal1 ;
  RECT 283.120 0.000 286.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal3 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal2 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal1 ;
  RECT 274.440 0.000 277.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 265.760 0.000 269.300 1.120 ;
  LAYER metal3 ;
  RECT 265.760 0.000 269.300 1.120 ;
  LAYER metal2 ;
  RECT 265.760 0.000 269.300 1.120 ;
  LAYER metal1 ;
  RECT 265.760 0.000 269.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal3 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal2 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal1 ;
  RECT 253.360 0.000 256.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 231.040 0.000 234.580 1.120 ;
  LAYER metal3 ;
  RECT 231.040 0.000 234.580 1.120 ;
  LAYER metal2 ;
  RECT 231.040 0.000 234.580 1.120 ;
  LAYER metal1 ;
  RECT 231.040 0.000 234.580 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 222.360 0.000 225.900 1.120 ;
  LAYER metal3 ;
  RECT 222.360 0.000 225.900 1.120 ;
  LAYER metal2 ;
  RECT 222.360 0.000 225.900 1.120 ;
  LAYER metal1 ;
  RECT 222.360 0.000 225.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 178.960 0.000 182.500 1.120 ;
  LAYER metal3 ;
  RECT 178.960 0.000 182.500 1.120 ;
  LAYER metal2 ;
  RECT 178.960 0.000 182.500 1.120 ;
  LAYER metal1 ;
  RECT 178.960 0.000 182.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 170.280 0.000 173.820 1.120 ;
  LAYER metal3 ;
  RECT 170.280 0.000 173.820 1.120 ;
  LAYER metal2 ;
  RECT 170.280 0.000 173.820 1.120 ;
  LAYER metal1 ;
  RECT 170.280 0.000 173.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 161.600 0.000 165.140 1.120 ;
  LAYER metal3 ;
  RECT 161.600 0.000 165.140 1.120 ;
  LAYER metal2 ;
  RECT 161.600 0.000 165.140 1.120 ;
  LAYER metal1 ;
  RECT 161.600 0.000 165.140 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 152.920 0.000 156.460 1.120 ;
  LAYER metal3 ;
  RECT 152.920 0.000 156.460 1.120 ;
  LAYER metal2 ;
  RECT 152.920 0.000 156.460 1.120 ;
  LAYER metal1 ;
  RECT 152.920 0.000 156.460 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 118.200 0.000 121.740 1.120 ;
  LAYER metal3 ;
  RECT 118.200 0.000 121.740 1.120 ;
  LAYER metal2 ;
  RECT 118.200 0.000 121.740 1.120 ;
  LAYER metal1 ;
  RECT 118.200 0.000 121.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 74.800 0.000 78.340 1.120 ;
  LAYER metal3 ;
  RECT 74.800 0.000 78.340 1.120 ;
  LAYER metal2 ;
  RECT 74.800 0.000 78.340 1.120 ;
  LAYER metal1 ;
  RECT 74.800 0.000 78.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 66.120 0.000 69.660 1.120 ;
  LAYER metal3 ;
  RECT 66.120 0.000 69.660 1.120 ;
  LAYER metal2 ;
  RECT 66.120 0.000 69.660 1.120 ;
  LAYER metal1 ;
  RECT 66.120 0.000 69.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER metal3 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER metal2 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER metal1 ;
  RECT 57.440 0.000 60.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER metal3 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER metal2 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER metal1 ;
  RECT 48.760 0.000 52.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER metal3 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER metal2 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER metal1 ;
  RECT 40.080 0.000 43.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN DO[31]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1819.760 0.000 1820.880 1.120 ;
  LAYER metal3 ;
  RECT 1819.760 0.000 1820.880 1.120 ;
  LAYER metal2 ;
  RECT 1819.760 0.000 1820.880 1.120 ;
  LAYER metal1 ;
  RECT 1819.760 0.000 1820.880 1.120 ;
 END
END DO[31]
PIN DI[31]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1811.700 0.000 1812.820 1.120 ;
  LAYER metal3 ;
  RECT 1811.700 0.000 1812.820 1.120 ;
  LAYER metal2 ;
  RECT 1811.700 0.000 1812.820 1.120 ;
  LAYER metal1 ;
  RECT 1811.700 0.000 1812.820 1.120 ;
 END
END DI[31]
PIN DO[30]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1806.740 0.000 1807.860 1.120 ;
  LAYER metal3 ;
  RECT 1806.740 0.000 1807.860 1.120 ;
  LAYER metal2 ;
  RECT 1806.740 0.000 1807.860 1.120 ;
  LAYER metal1 ;
  RECT 1806.740 0.000 1807.860 1.120 ;
 END
END DO[30]
PIN DI[30]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1798.060 0.000 1799.180 1.120 ;
  LAYER metal3 ;
  RECT 1798.060 0.000 1799.180 1.120 ;
  LAYER metal2 ;
  RECT 1798.060 0.000 1799.180 1.120 ;
  LAYER metal1 ;
  RECT 1798.060 0.000 1799.180 1.120 ;
 END
END DI[30]
PIN DO[29]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1706.920 0.000 1708.040 1.120 ;
  LAYER metal3 ;
  RECT 1706.920 0.000 1708.040 1.120 ;
  LAYER metal2 ;
  RECT 1706.920 0.000 1708.040 1.120 ;
  LAYER metal1 ;
  RECT 1706.920 0.000 1708.040 1.120 ;
 END
END DO[29]
PIN DI[29]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1698.860 0.000 1699.980 1.120 ;
  LAYER metal3 ;
  RECT 1698.860 0.000 1699.980 1.120 ;
  LAYER metal2 ;
  RECT 1698.860 0.000 1699.980 1.120 ;
  LAYER metal1 ;
  RECT 1698.860 0.000 1699.980 1.120 ;
 END
END DI[29]
PIN DO[28]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1693.900 0.000 1695.020 1.120 ;
  LAYER metal3 ;
  RECT 1693.900 0.000 1695.020 1.120 ;
  LAYER metal2 ;
  RECT 1693.900 0.000 1695.020 1.120 ;
  LAYER metal1 ;
  RECT 1693.900 0.000 1695.020 1.120 ;
 END
END DO[28]
PIN DI[28]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1685.220 0.000 1686.340 1.120 ;
  LAYER metal3 ;
  RECT 1685.220 0.000 1686.340 1.120 ;
  LAYER metal2 ;
  RECT 1685.220 0.000 1686.340 1.120 ;
  LAYER metal1 ;
  RECT 1685.220 0.000 1686.340 1.120 ;
 END
END DI[28]
PIN DO[27]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1594.080 0.000 1595.200 1.120 ;
  LAYER metal3 ;
  RECT 1594.080 0.000 1595.200 1.120 ;
  LAYER metal2 ;
  RECT 1594.080 0.000 1595.200 1.120 ;
  LAYER metal1 ;
  RECT 1594.080 0.000 1595.200 1.120 ;
 END
END DO[27]
PIN DI[27]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal3 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal2 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal1 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
 END
END DI[27]
PIN DO[26]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1580.440 0.000 1581.560 1.120 ;
  LAYER metal3 ;
  RECT 1580.440 0.000 1581.560 1.120 ;
  LAYER metal2 ;
  RECT 1580.440 0.000 1581.560 1.120 ;
  LAYER metal1 ;
  RECT 1580.440 0.000 1581.560 1.120 ;
 END
END DO[26]
PIN DI[26]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1572.380 0.000 1573.500 1.120 ;
  LAYER metal3 ;
  RECT 1572.380 0.000 1573.500 1.120 ;
  LAYER metal2 ;
  RECT 1572.380 0.000 1573.500 1.120 ;
  LAYER metal1 ;
  RECT 1572.380 0.000 1573.500 1.120 ;
 END
END DI[26]
PIN DO[25]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1480.620 0.000 1481.740 1.120 ;
  LAYER metal3 ;
  RECT 1480.620 0.000 1481.740 1.120 ;
  LAYER metal2 ;
  RECT 1480.620 0.000 1481.740 1.120 ;
  LAYER metal1 ;
  RECT 1480.620 0.000 1481.740 1.120 ;
 END
END DO[25]
PIN DI[25]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1472.560 0.000 1473.680 1.120 ;
  LAYER metal3 ;
  RECT 1472.560 0.000 1473.680 1.120 ;
  LAYER metal2 ;
  RECT 1472.560 0.000 1473.680 1.120 ;
  LAYER metal1 ;
  RECT 1472.560 0.000 1473.680 1.120 ;
 END
END DI[25]
PIN DO[24]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1467.600 0.000 1468.720 1.120 ;
  LAYER metal3 ;
  RECT 1467.600 0.000 1468.720 1.120 ;
  LAYER metal2 ;
  RECT 1467.600 0.000 1468.720 1.120 ;
  LAYER metal1 ;
  RECT 1467.600 0.000 1468.720 1.120 ;
 END
END DO[24]
PIN DI[24]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1458.920 0.000 1460.040 1.120 ;
  LAYER metal3 ;
  RECT 1458.920 0.000 1460.040 1.120 ;
  LAYER metal2 ;
  RECT 1458.920 0.000 1460.040 1.120 ;
  LAYER metal1 ;
  RECT 1458.920 0.000 1460.040 1.120 ;
 END
END DI[24]
PIN DO[23]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1367.780 0.000 1368.900 1.120 ;
  LAYER metal3 ;
  RECT 1367.780 0.000 1368.900 1.120 ;
  LAYER metal2 ;
  RECT 1367.780 0.000 1368.900 1.120 ;
  LAYER metal1 ;
  RECT 1367.780 0.000 1368.900 1.120 ;
 END
END DO[23]
PIN DI[23]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1359.720 0.000 1360.840 1.120 ;
  LAYER metal3 ;
  RECT 1359.720 0.000 1360.840 1.120 ;
  LAYER metal2 ;
  RECT 1359.720 0.000 1360.840 1.120 ;
  LAYER metal1 ;
  RECT 1359.720 0.000 1360.840 1.120 ;
 END
END DI[23]
PIN DO[22]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1354.760 0.000 1355.880 1.120 ;
  LAYER metal3 ;
  RECT 1354.760 0.000 1355.880 1.120 ;
  LAYER metal2 ;
  RECT 1354.760 0.000 1355.880 1.120 ;
  LAYER metal1 ;
  RECT 1354.760 0.000 1355.880 1.120 ;
 END
END DO[22]
PIN DI[22]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1346.080 0.000 1347.200 1.120 ;
  LAYER metal3 ;
  RECT 1346.080 0.000 1347.200 1.120 ;
  LAYER metal2 ;
  RECT 1346.080 0.000 1347.200 1.120 ;
  LAYER metal1 ;
  RECT 1346.080 0.000 1347.200 1.120 ;
 END
END DI[22]
PIN DO[21]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1254.940 0.000 1256.060 1.120 ;
  LAYER metal3 ;
  RECT 1254.940 0.000 1256.060 1.120 ;
  LAYER metal2 ;
  RECT 1254.940 0.000 1256.060 1.120 ;
  LAYER metal1 ;
  RECT 1254.940 0.000 1256.060 1.120 ;
 END
END DO[21]
PIN DI[21]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1246.260 0.000 1247.380 1.120 ;
  LAYER metal3 ;
  RECT 1246.260 0.000 1247.380 1.120 ;
  LAYER metal2 ;
  RECT 1246.260 0.000 1247.380 1.120 ;
  LAYER metal1 ;
  RECT 1246.260 0.000 1247.380 1.120 ;
 END
END DI[21]
PIN DO[20]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1241.300 0.000 1242.420 1.120 ;
  LAYER metal3 ;
  RECT 1241.300 0.000 1242.420 1.120 ;
  LAYER metal2 ;
  RECT 1241.300 0.000 1242.420 1.120 ;
  LAYER metal1 ;
  RECT 1241.300 0.000 1242.420 1.120 ;
 END
END DO[20]
PIN DI[20]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1233.240 0.000 1234.360 1.120 ;
  LAYER metal3 ;
  RECT 1233.240 0.000 1234.360 1.120 ;
  LAYER metal2 ;
  RECT 1233.240 0.000 1234.360 1.120 ;
  LAYER metal1 ;
  RECT 1233.240 0.000 1234.360 1.120 ;
 END
END DI[20]
PIN DO[19]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal3 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal2 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal1 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
 END
END DO[19]
PIN DI[19]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1133.420 0.000 1134.540 1.120 ;
  LAYER metal3 ;
  RECT 1133.420 0.000 1134.540 1.120 ;
  LAYER metal2 ;
  RECT 1133.420 0.000 1134.540 1.120 ;
  LAYER metal1 ;
  RECT 1133.420 0.000 1134.540 1.120 ;
 END
END DI[19]
PIN DO[18]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal3 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal2 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal1 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
 END
END DO[18]
PIN DI[18]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1119.780 0.000 1120.900 1.120 ;
  LAYER metal3 ;
  RECT 1119.780 0.000 1120.900 1.120 ;
  LAYER metal2 ;
  RECT 1119.780 0.000 1120.900 1.120 ;
  LAYER metal1 ;
  RECT 1119.780 0.000 1120.900 1.120 ;
 END
END DI[18]
PIN DO[17]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1028.640 0.000 1029.760 1.120 ;
  LAYER metal3 ;
  RECT 1028.640 0.000 1029.760 1.120 ;
  LAYER metal2 ;
  RECT 1028.640 0.000 1029.760 1.120 ;
  LAYER metal1 ;
  RECT 1028.640 0.000 1029.760 1.120 ;
 END
END DO[17]
PIN DI[17]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal3 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal2 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal1 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
 END
END DI[17]
PIN DO[16]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1015.620 0.000 1016.740 1.120 ;
  LAYER metal3 ;
  RECT 1015.620 0.000 1016.740 1.120 ;
  LAYER metal2 ;
  RECT 1015.620 0.000 1016.740 1.120 ;
  LAYER metal1 ;
  RECT 1015.620 0.000 1016.740 1.120 ;
 END
END DO[16]
PIN DI[16]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1006.940 0.000 1008.060 1.120 ;
  LAYER metal3 ;
  RECT 1006.940 0.000 1008.060 1.120 ;
  LAYER metal2 ;
  RECT 1006.940 0.000 1008.060 1.120 ;
  LAYER metal1 ;
  RECT 1006.940 0.000 1008.060 1.120 ;
 END
END DI[16]
PIN A[1]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 1001.360 0.000 1002.480 1.120 ;
  LAYER metal3 ;
  RECT 1001.360 0.000 1002.480 1.120 ;
  LAYER metal2 ;
  RECT 1001.360 0.000 1002.480 1.120 ;
  LAYER metal1 ;
  RECT 1001.360 0.000 1002.480 1.120 ;
 END
END A[1]
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 999.500 0.000 1000.620 1.120 ;
  LAYER metal3 ;
  RECT 999.500 0.000 1000.620 1.120 ;
  LAYER metal2 ;
  RECT 999.500 0.000 1000.620 1.120 ;
  LAYER metal1 ;
  RECT 999.500 0.000 1000.620 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER metal4 ;
  RECT 994.540 0.000 995.660 1.120 ;
  LAYER metal3 ;
  RECT 994.540 0.000 995.660 1.120 ;
  LAYER metal2 ;
  RECT 994.540 0.000 995.660 1.120 ;
  LAYER metal1 ;
  RECT 994.540 0.000 995.660 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER metal4 ;
  RECT 992.680 0.000 993.800 1.120 ;
  LAYER metal3 ;
  RECT 992.680 0.000 993.800 1.120 ;
  LAYER metal2 ;
  RECT 992.680 0.000 993.800 1.120 ;
  LAYER metal1 ;
  RECT 992.680 0.000 993.800 1.120 ;
 END
END CS
PIN A[3]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 990.820 0.000 991.940 1.120 ;
  LAYER metal3 ;
  RECT 990.820 0.000 991.940 1.120 ;
  LAYER metal2 ;
  RECT 990.820 0.000 991.940 1.120 ;
  LAYER metal1 ;
  RECT 990.820 0.000 991.940 1.120 ;
 END
END A[3]
PIN A[4]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 984.000 0.000 985.120 1.120 ;
  LAYER metal3 ;
  RECT 984.000 0.000 985.120 1.120 ;
  LAYER metal2 ;
  RECT 984.000 0.000 985.120 1.120 ;
  LAYER metal1 ;
  RECT 984.000 0.000 985.120 1.120 ;
 END
END A[4]
PIN A[2]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 970.980 0.000 972.100 1.120 ;
  LAYER metal3 ;
  RECT 970.980 0.000 972.100 1.120 ;
  LAYER metal2 ;
  RECT 970.980 0.000 972.100 1.120 ;
  LAYER metal1 ;
  RECT 970.980 0.000 972.100 1.120 ;
 END
END A[2]
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER metal4 ;
  RECT 968.500 0.000 969.620 1.120 ;
  LAYER metal3 ;
  RECT 968.500 0.000 969.620 1.120 ;
  LAYER metal2 ;
  RECT 968.500 0.000 969.620 1.120 ;
  LAYER metal1 ;
  RECT 968.500 0.000 969.620 1.120 ;
 END
END CK
PIN A[0]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 966.020 0.000 967.140 1.120 ;
  LAYER metal3 ;
  RECT 966.020 0.000 967.140 1.120 ;
  LAYER metal2 ;
  RECT 966.020 0.000 967.140 1.120 ;
  LAYER metal1 ;
  RECT 966.020 0.000 967.140 1.120 ;
 END
END A[0]
PIN A[5]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 961.680 0.000 962.800 1.120 ;
  LAYER metal3 ;
  RECT 961.680 0.000 962.800 1.120 ;
  LAYER metal2 ;
  RECT 961.680 0.000 962.800 1.120 ;
  LAYER metal1 ;
  RECT 961.680 0.000 962.800 1.120 ;
 END
END A[5]
PIN A[6]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 954.240 0.000 955.360 1.120 ;
  LAYER metal3 ;
  RECT 954.240 0.000 955.360 1.120 ;
  LAYER metal2 ;
  RECT 954.240 0.000 955.360 1.120 ;
  LAYER metal1 ;
  RECT 954.240 0.000 955.360 1.120 ;
 END
END A[6]
PIN A[7]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 951.140 0.000 952.260 1.120 ;
  LAYER metal3 ;
  RECT 951.140 0.000 952.260 1.120 ;
  LAYER metal2 ;
  RECT 951.140 0.000 952.260 1.120 ;
  LAYER metal1 ;
  RECT 951.140 0.000 952.260 1.120 ;
 END
END A[7]
PIN A[8]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 943.700 0.000 944.820 1.120 ;
  LAYER metal3 ;
  RECT 943.700 0.000 944.820 1.120 ;
  LAYER metal2 ;
  RECT 943.700 0.000 944.820 1.120 ;
  LAYER metal1 ;
  RECT 943.700 0.000 944.820 1.120 ;
 END
END A[8]
PIN A[9]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 940.600 0.000 941.720 1.120 ;
  LAYER metal3 ;
  RECT 940.600 0.000 941.720 1.120 ;
  LAYER metal2 ;
  RECT 940.600 0.000 941.720 1.120 ;
  LAYER metal1 ;
  RECT 940.600 0.000 941.720 1.120 ;
 END
END A[9]
PIN A[10]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 933.160 0.000 934.280 1.120 ;
  LAYER metal3 ;
  RECT 933.160 0.000 934.280 1.120 ;
  LAYER metal2 ;
  RECT 933.160 0.000 934.280 1.120 ;
  LAYER metal1 ;
  RECT 933.160 0.000 934.280 1.120 ;
 END
END A[10]
PIN A[11]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 930.060 0.000 931.180 1.120 ;
  LAYER metal3 ;
  RECT 930.060 0.000 931.180 1.120 ;
  LAYER metal2 ;
  RECT 930.060 0.000 931.180 1.120 ;
  LAYER metal1 ;
  RECT 930.060 0.000 931.180 1.120 ;
 END
END A[11]
PIN A[12]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 922.000 0.000 923.120 1.120 ;
  LAYER metal3 ;
  RECT 922.000 0.000 923.120 1.120 ;
  LAYER metal2 ;
  RECT 922.000 0.000 923.120 1.120 ;
  LAYER metal1 ;
  RECT 922.000 0.000 923.120 1.120 ;
 END
END A[12]
PIN A[13]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 919.520 0.000 920.640 1.120 ;
  LAYER metal3 ;
  RECT 919.520 0.000 920.640 1.120 ;
  LAYER metal2 ;
  RECT 919.520 0.000 920.640 1.120 ;
  LAYER metal1 ;
  RECT 919.520 0.000 920.640 1.120 ;
 END
END A[13]
PIN DO[15]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 824.660 0.000 825.780 1.120 ;
  LAYER metal3 ;
  RECT 824.660 0.000 825.780 1.120 ;
  LAYER metal2 ;
  RECT 824.660 0.000 825.780 1.120 ;
  LAYER metal1 ;
  RECT 824.660 0.000 825.780 1.120 ;
 END
END DO[15]
PIN DI[15]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 815.980 0.000 817.100 1.120 ;
  LAYER metal3 ;
  RECT 815.980 0.000 817.100 1.120 ;
  LAYER metal2 ;
  RECT 815.980 0.000 817.100 1.120 ;
  LAYER metal1 ;
  RECT 815.980 0.000 817.100 1.120 ;
 END
END DI[15]
PIN DO[14]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 811.640 0.000 812.760 1.120 ;
  LAYER metal3 ;
  RECT 811.640 0.000 812.760 1.120 ;
  LAYER metal2 ;
  RECT 811.640 0.000 812.760 1.120 ;
  LAYER metal1 ;
  RECT 811.640 0.000 812.760 1.120 ;
 END
END DO[14]
PIN DI[14]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 802.960 0.000 804.080 1.120 ;
  LAYER metal3 ;
  RECT 802.960 0.000 804.080 1.120 ;
  LAYER metal2 ;
  RECT 802.960 0.000 804.080 1.120 ;
  LAYER metal1 ;
  RECT 802.960 0.000 804.080 1.120 ;
 END
END DI[14]
PIN DO[13]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal3 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal2 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal1 ;
  RECT 711.820 0.000 712.940 1.120 ;
 END
END DO[13]
PIN DI[13]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 703.140 0.000 704.260 1.120 ;
  LAYER metal3 ;
  RECT 703.140 0.000 704.260 1.120 ;
  LAYER metal2 ;
  RECT 703.140 0.000 704.260 1.120 ;
  LAYER metal1 ;
  RECT 703.140 0.000 704.260 1.120 ;
 END
END DI[13]
PIN DO[12]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal3 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal2 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal1 ;
  RECT 698.180 0.000 699.300 1.120 ;
 END
END DO[12]
PIN DI[12]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 690.120 0.000 691.240 1.120 ;
  LAYER metal3 ;
  RECT 690.120 0.000 691.240 1.120 ;
  LAYER metal2 ;
  RECT 690.120 0.000 691.240 1.120 ;
  LAYER metal1 ;
  RECT 690.120 0.000 691.240 1.120 ;
 END
END DI[12]
PIN DO[11]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER metal3 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER metal2 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER metal1 ;
  RECT 598.360 0.000 599.480 1.120 ;
 END
END DO[11]
PIN DI[11]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER metal3 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER metal2 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER metal1 ;
  RECT 590.300 0.000 591.420 1.120 ;
 END
END DI[11]
PIN DO[10]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER metal3 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER metal2 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER metal1 ;
  RECT 585.340 0.000 586.460 1.120 ;
 END
END DO[10]
PIN DI[10]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER metal3 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER metal2 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER metal1 ;
  RECT 576.660 0.000 577.780 1.120 ;
 END
END DI[10]
PIN DO[9]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER metal3 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER metal2 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER metal1 ;
  RECT 485.520 0.000 486.640 1.120 ;
 END
END DO[9]
PIN DI[9]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER metal3 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER metal2 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER metal1 ;
  RECT 476.840 0.000 477.960 1.120 ;
 END
END DI[9]
PIN DO[8]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER metal3 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER metal2 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER metal1 ;
  RECT 472.500 0.000 473.620 1.120 ;
 END
END DO[8]
PIN DI[8]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER metal3 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER metal2 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER metal1 ;
  RECT 463.820 0.000 464.940 1.120 ;
 END
END DI[8]
PIN DO[7]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER metal3 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER metal2 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER metal1 ;
  RECT 372.680 0.000 373.800 1.120 ;
 END
END DO[7]
PIN DI[7]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER metal3 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER metal2 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER metal1 ;
  RECT 364.000 0.000 365.120 1.120 ;
 END
END DI[7]
PIN DO[6]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal3 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal2 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal1 ;
  RECT 359.040 0.000 360.160 1.120 ;
 END
END DO[6]
PIN DI[6]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER metal3 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER metal2 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER metal1 ;
  RECT 350.980 0.000 352.100 1.120 ;
 END
END DI[6]
PIN DO[5]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DO[5]
PIN DI[5]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal3 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal2 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal1 ;
  RECT 251.160 0.000 252.280 1.120 ;
 END
END DI[5]
PIN DO[4]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal3 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal2 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal1 ;
  RECT 246.200 0.000 247.320 1.120 ;
 END
END DO[4]
PIN DI[4]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal3 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal2 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal1 ;
  RECT 237.520 0.000 238.640 1.120 ;
 END
END DI[4]
PIN DO[3]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO[3]
PIN DI[3]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI[3]
PIN DO[2]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO[2]
PIN DI[2]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI[2]
PIN DO[1]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO[1]
PIN DI[1]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI[1]
PIN DO[0]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO[0]
PIN DI[0]
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI[0]
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 1920.140 1391.600 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 1920.140 1391.600 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 1920.140 1391.600 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 1920.140 1391.600 ;
  LAYER via ;
  RECT 0.000 0.140 1920.140 1391.600 ;
  LAYER via2 ;
  RECT 0.000 0.140 1920.140 1391.600 ;
  LAYER via3 ;
  RECT 0.000 0.140 1920.140 1391.600 ;
END
END SRAM
END LIBRARY



